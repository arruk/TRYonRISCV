TORVS/torvs9C.sv