TORVS/torvs7C.sv