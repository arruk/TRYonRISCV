//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.10.03 Education
//Part Number: GW5A-LV25MG121NC1/I0
//Device: GW5A-25
//Device Version: A
//Created Time: Wed Jan  8 20:44:32 2025

module Gowin_DPB (douta, doutb, clka, ocea, cea, reseta, wrea, clkb, oceb, ceb, resetb, wreb, ada, dina, adb, dinb, byte_ena, byte_enb);

output [31:0] douta;
output [31:0] doutb;
input clka;
input ocea;
input cea;
input reseta;
input wrea;
input clkb;
input oceb;
input ceb;
input resetb;
input wreb;
input [13:0] ada;
input [31:0] dina;
input [13:0] adb;
input [31:0] dinb;
input [3:0] byte_ena;
input [3:0] byte_enb;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire lut_f_10;
wire lut_f_11;
wire lut_f_12;
wire lut_f_13;
wire lut_f_14;
wire lut_f_15;
wire lut_f_16;
wire lut_f_17;
wire lut_f_18;
wire lut_f_19;
wire lut_f_20;
wire lut_f_21;
wire lut_f_22;
wire lut_f_23;
wire lut_f_24;
wire lut_f_25;
wire lut_f_26;
wire lut_f_27;
wire lut_f_28;
wire lut_f_29;
wire lut_f_30;
wire lut_f_31;
wire [15:0] dpb_inst_0_douta;
wire [15:0] dpb_inst_0_doutb;
wire [15:0] dpb_inst_1_douta;
wire [15:0] dpb_inst_1_doutb;
wire [15:0] dpb_inst_2_douta;
wire [15:0] dpb_inst_2_doutb;
wire [15:0] dpb_inst_3_douta;
wire [15:0] dpb_inst_3_doutb;
wire [15:0] dpb_inst_4_douta;
wire [15:0] dpb_inst_4_doutb;
wire [15:0] dpb_inst_5_douta;
wire [15:0] dpb_inst_5_doutb;
wire [15:0] dpb_inst_6_douta;
wire [15:0] dpb_inst_6_doutb;
wire [15:0] dpb_inst_7_douta;
wire [15:0] dpb_inst_7_doutb;
wire [15:0] dpb_inst_8_douta;
wire [15:0] dpb_inst_8_doutb;
wire [15:0] dpb_inst_9_douta;
wire [15:0] dpb_inst_9_doutb;
wire [15:0] dpb_inst_10_douta;
wire [15:0] dpb_inst_10_doutb;
wire [15:0] dpb_inst_11_douta;
wire [15:0] dpb_inst_11_doutb;
wire [15:0] dpb_inst_12_douta;
wire [15:0] dpb_inst_12_doutb;
wire [15:0] dpb_inst_13_douta;
wire [15:0] dpb_inst_13_doutb;
wire [15:0] dpb_inst_14_douta;
wire [15:0] dpb_inst_14_doutb;
wire [15:0] dpb_inst_15_douta;
wire [15:0] dpb_inst_15_doutb;
wire [31:16] dpb_inst_16_douta;
wire [31:16] dpb_inst_16_doutb;
wire [31:16] dpb_inst_17_douta;
wire [31:16] dpb_inst_17_doutb;
wire [31:16] dpb_inst_18_douta;
wire [31:16] dpb_inst_18_doutb;
wire [31:16] dpb_inst_19_douta;
wire [31:16] dpb_inst_19_doutb;
wire [31:16] dpb_inst_20_douta;
wire [31:16] dpb_inst_20_doutb;
wire [31:16] dpb_inst_21_douta;
wire [31:16] dpb_inst_21_doutb;
wire [31:16] dpb_inst_22_douta;
wire [31:16] dpb_inst_22_doutb;
wire [31:16] dpb_inst_23_douta;
wire [31:16] dpb_inst_23_doutb;
wire [31:16] dpb_inst_24_douta;
wire [31:16] dpb_inst_24_doutb;
wire [31:16] dpb_inst_25_douta;
wire [31:16] dpb_inst_25_doutb;
wire [31:16] dpb_inst_26_douta;
wire [31:16] dpb_inst_26_doutb;
wire [31:16] dpb_inst_27_douta;
wire [31:16] dpb_inst_27_doutb;
wire [31:16] dpb_inst_28_douta;
wire [31:16] dpb_inst_28_doutb;
wire [31:16] dpb_inst_29_douta;
wire [31:16] dpb_inst_29_doutb;
wire [31:16] dpb_inst_30_douta;
wire [31:16] dpb_inst_30_doutb;
wire [31:16] dpb_inst_31_douta;
wire [31:16] dpb_inst_31_doutb;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire dff_q_4;
wire dff_q_5;
wire dff_q_6;
wire dff_q_7;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;
wire mux_o_6;
wire mux_o_7;
wire mux_o_8;
wire mux_o_9;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_13;
wire mux_o_15;
wire mux_o_16;
wire mux_o_17;
wire mux_o_18;
wire mux_o_19;
wire mux_o_20;
wire mux_o_21;
wire mux_o_22;
wire mux_o_23;
wire mux_o_24;
wire mux_o_25;
wire mux_o_26;
wire mux_o_27;
wire mux_o_28;
wire mux_o_30;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_34;
wire mux_o_35;
wire mux_o_36;
wire mux_o_37;
wire mux_o_38;
wire mux_o_39;
wire mux_o_40;
wire mux_o_41;
wire mux_o_42;
wire mux_o_43;
wire mux_o_45;
wire mux_o_46;
wire mux_o_47;
wire mux_o_48;
wire mux_o_49;
wire mux_o_50;
wire mux_o_51;
wire mux_o_52;
wire mux_o_53;
wire mux_o_54;
wire mux_o_55;
wire mux_o_56;
wire mux_o_57;
wire mux_o_58;
wire mux_o_60;
wire mux_o_61;
wire mux_o_62;
wire mux_o_63;
wire mux_o_64;
wire mux_o_65;
wire mux_o_66;
wire mux_o_67;
wire mux_o_68;
wire mux_o_69;
wire mux_o_70;
wire mux_o_71;
wire mux_o_72;
wire mux_o_73;
wire mux_o_75;
wire mux_o_76;
wire mux_o_77;
wire mux_o_78;
wire mux_o_79;
wire mux_o_80;
wire mux_o_81;
wire mux_o_82;
wire mux_o_83;
wire mux_o_84;
wire mux_o_85;
wire mux_o_86;
wire mux_o_87;
wire mux_o_88;
wire mux_o_90;
wire mux_o_91;
wire mux_o_92;
wire mux_o_93;
wire mux_o_94;
wire mux_o_95;
wire mux_o_96;
wire mux_o_97;
wire mux_o_98;
wire mux_o_99;
wire mux_o_100;
wire mux_o_101;
wire mux_o_102;
wire mux_o_103;
wire mux_o_105;
wire mux_o_106;
wire mux_o_107;
wire mux_o_108;
wire mux_o_109;
wire mux_o_110;
wire mux_o_111;
wire mux_o_112;
wire mux_o_113;
wire mux_o_114;
wire mux_o_115;
wire mux_o_116;
wire mux_o_117;
wire mux_o_118;
wire mux_o_120;
wire mux_o_121;
wire mux_o_122;
wire mux_o_123;
wire mux_o_124;
wire mux_o_125;
wire mux_o_126;
wire mux_o_127;
wire mux_o_128;
wire mux_o_129;
wire mux_o_130;
wire mux_o_131;
wire mux_o_132;
wire mux_o_133;
wire mux_o_135;
wire mux_o_136;
wire mux_o_137;
wire mux_o_138;
wire mux_o_139;
wire mux_o_140;
wire mux_o_141;
wire mux_o_142;
wire mux_o_143;
wire mux_o_144;
wire mux_o_145;
wire mux_o_146;
wire mux_o_147;
wire mux_o_148;
wire mux_o_150;
wire mux_o_151;
wire mux_o_152;
wire mux_o_153;
wire mux_o_154;
wire mux_o_155;
wire mux_o_156;
wire mux_o_157;
wire mux_o_158;
wire mux_o_159;
wire mux_o_160;
wire mux_o_161;
wire mux_o_162;
wire mux_o_163;
wire mux_o_165;
wire mux_o_166;
wire mux_o_167;
wire mux_o_168;
wire mux_o_169;
wire mux_o_170;
wire mux_o_171;
wire mux_o_172;
wire mux_o_173;
wire mux_o_174;
wire mux_o_175;
wire mux_o_176;
wire mux_o_177;
wire mux_o_178;
wire mux_o_180;
wire mux_o_181;
wire mux_o_182;
wire mux_o_183;
wire mux_o_184;
wire mux_o_185;
wire mux_o_186;
wire mux_o_187;
wire mux_o_188;
wire mux_o_189;
wire mux_o_190;
wire mux_o_191;
wire mux_o_192;
wire mux_o_193;
wire mux_o_195;
wire mux_o_196;
wire mux_o_197;
wire mux_o_198;
wire mux_o_199;
wire mux_o_200;
wire mux_o_201;
wire mux_o_202;
wire mux_o_203;
wire mux_o_204;
wire mux_o_205;
wire mux_o_206;
wire mux_o_207;
wire mux_o_208;
wire mux_o_210;
wire mux_o_211;
wire mux_o_212;
wire mux_o_213;
wire mux_o_214;
wire mux_o_215;
wire mux_o_216;
wire mux_o_217;
wire mux_o_218;
wire mux_o_219;
wire mux_o_220;
wire mux_o_221;
wire mux_o_222;
wire mux_o_223;
wire mux_o_225;
wire mux_o_226;
wire mux_o_227;
wire mux_o_228;
wire mux_o_229;
wire mux_o_230;
wire mux_o_231;
wire mux_o_232;
wire mux_o_233;
wire mux_o_234;
wire mux_o_235;
wire mux_o_236;
wire mux_o_237;
wire mux_o_238;
wire mux_o_240;
wire mux_o_241;
wire mux_o_242;
wire mux_o_243;
wire mux_o_244;
wire mux_o_245;
wire mux_o_246;
wire mux_o_247;
wire mux_o_248;
wire mux_o_249;
wire mux_o_250;
wire mux_o_251;
wire mux_o_252;
wire mux_o_253;
wire mux_o_255;
wire mux_o_256;
wire mux_o_257;
wire mux_o_258;
wire mux_o_259;
wire mux_o_260;
wire mux_o_261;
wire mux_o_262;
wire mux_o_263;
wire mux_o_264;
wire mux_o_265;
wire mux_o_266;
wire mux_o_267;
wire mux_o_268;
wire mux_o_270;
wire mux_o_271;
wire mux_o_272;
wire mux_o_273;
wire mux_o_274;
wire mux_o_275;
wire mux_o_276;
wire mux_o_277;
wire mux_o_278;
wire mux_o_279;
wire mux_o_280;
wire mux_o_281;
wire mux_o_282;
wire mux_o_283;
wire mux_o_285;
wire mux_o_286;
wire mux_o_287;
wire mux_o_288;
wire mux_o_289;
wire mux_o_290;
wire mux_o_291;
wire mux_o_292;
wire mux_o_293;
wire mux_o_294;
wire mux_o_295;
wire mux_o_296;
wire mux_o_297;
wire mux_o_298;
wire mux_o_300;
wire mux_o_301;
wire mux_o_302;
wire mux_o_303;
wire mux_o_304;
wire mux_o_305;
wire mux_o_306;
wire mux_o_307;
wire mux_o_308;
wire mux_o_309;
wire mux_o_310;
wire mux_o_311;
wire mux_o_312;
wire mux_o_313;
wire mux_o_315;
wire mux_o_316;
wire mux_o_317;
wire mux_o_318;
wire mux_o_319;
wire mux_o_320;
wire mux_o_321;
wire mux_o_322;
wire mux_o_323;
wire mux_o_324;
wire mux_o_325;
wire mux_o_326;
wire mux_o_327;
wire mux_o_328;
wire mux_o_330;
wire mux_o_331;
wire mux_o_332;
wire mux_o_333;
wire mux_o_334;
wire mux_o_335;
wire mux_o_336;
wire mux_o_337;
wire mux_o_338;
wire mux_o_339;
wire mux_o_340;
wire mux_o_341;
wire mux_o_342;
wire mux_o_343;
wire mux_o_345;
wire mux_o_346;
wire mux_o_347;
wire mux_o_348;
wire mux_o_349;
wire mux_o_350;
wire mux_o_351;
wire mux_o_352;
wire mux_o_353;
wire mux_o_354;
wire mux_o_355;
wire mux_o_356;
wire mux_o_357;
wire mux_o_358;
wire mux_o_360;
wire mux_o_361;
wire mux_o_362;
wire mux_o_363;
wire mux_o_364;
wire mux_o_365;
wire mux_o_366;
wire mux_o_367;
wire mux_o_368;
wire mux_o_369;
wire mux_o_370;
wire mux_o_371;
wire mux_o_372;
wire mux_o_373;
wire mux_o_375;
wire mux_o_376;
wire mux_o_377;
wire mux_o_378;
wire mux_o_379;
wire mux_o_380;
wire mux_o_381;
wire mux_o_382;
wire mux_o_383;
wire mux_o_384;
wire mux_o_385;
wire mux_o_386;
wire mux_o_387;
wire mux_o_388;
wire mux_o_390;
wire mux_o_391;
wire mux_o_392;
wire mux_o_393;
wire mux_o_394;
wire mux_o_395;
wire mux_o_396;
wire mux_o_397;
wire mux_o_398;
wire mux_o_399;
wire mux_o_400;
wire mux_o_401;
wire mux_o_402;
wire mux_o_403;
wire mux_o_405;
wire mux_o_406;
wire mux_o_407;
wire mux_o_408;
wire mux_o_409;
wire mux_o_410;
wire mux_o_411;
wire mux_o_412;
wire mux_o_413;
wire mux_o_414;
wire mux_o_415;
wire mux_o_416;
wire mux_o_417;
wire mux_o_418;
wire mux_o_420;
wire mux_o_421;
wire mux_o_422;
wire mux_o_423;
wire mux_o_424;
wire mux_o_425;
wire mux_o_426;
wire mux_o_427;
wire mux_o_428;
wire mux_o_429;
wire mux_o_430;
wire mux_o_431;
wire mux_o_432;
wire mux_o_433;
wire mux_o_435;
wire mux_o_436;
wire mux_o_437;
wire mux_o_438;
wire mux_o_439;
wire mux_o_440;
wire mux_o_441;
wire mux_o_442;
wire mux_o_443;
wire mux_o_444;
wire mux_o_445;
wire mux_o_446;
wire mux_o_447;
wire mux_o_448;
wire mux_o_450;
wire mux_o_451;
wire mux_o_452;
wire mux_o_453;
wire mux_o_454;
wire mux_o_455;
wire mux_o_456;
wire mux_o_457;
wire mux_o_458;
wire mux_o_459;
wire mux_o_460;
wire mux_o_461;
wire mux_o_462;
wire mux_o_463;
wire mux_o_465;
wire mux_o_466;
wire mux_o_467;
wire mux_o_468;
wire mux_o_469;
wire mux_o_470;
wire mux_o_471;
wire mux_o_472;
wire mux_o_473;
wire mux_o_474;
wire mux_o_475;
wire mux_o_476;
wire mux_o_477;
wire mux_o_478;
wire mux_o_480;
wire mux_o_481;
wire mux_o_482;
wire mux_o_483;
wire mux_o_484;
wire mux_o_485;
wire mux_o_486;
wire mux_o_487;
wire mux_o_488;
wire mux_o_489;
wire mux_o_490;
wire mux_o_491;
wire mux_o_492;
wire mux_o_493;
wire mux_o_495;
wire mux_o_496;
wire mux_o_497;
wire mux_o_498;
wire mux_o_499;
wire mux_o_500;
wire mux_o_501;
wire mux_o_502;
wire mux_o_503;
wire mux_o_504;
wire mux_o_505;
wire mux_o_506;
wire mux_o_507;
wire mux_o_508;
wire mux_o_510;
wire mux_o_511;
wire mux_o_512;
wire mux_o_513;
wire mux_o_514;
wire mux_o_515;
wire mux_o_516;
wire mux_o_517;
wire mux_o_518;
wire mux_o_519;
wire mux_o_520;
wire mux_o_521;
wire mux_o_522;
wire mux_o_523;
wire mux_o_525;
wire mux_o_526;
wire mux_o_527;
wire mux_o_528;
wire mux_o_529;
wire mux_o_530;
wire mux_o_531;
wire mux_o_532;
wire mux_o_533;
wire mux_o_534;
wire mux_o_535;
wire mux_o_536;
wire mux_o_537;
wire mux_o_538;
wire mux_o_540;
wire mux_o_541;
wire mux_o_542;
wire mux_o_543;
wire mux_o_544;
wire mux_o_545;
wire mux_o_546;
wire mux_o_547;
wire mux_o_548;
wire mux_o_549;
wire mux_o_550;
wire mux_o_551;
wire mux_o_552;
wire mux_o_553;
wire mux_o_555;
wire mux_o_556;
wire mux_o_557;
wire mux_o_558;
wire mux_o_559;
wire mux_o_560;
wire mux_o_561;
wire mux_o_562;
wire mux_o_563;
wire mux_o_564;
wire mux_o_565;
wire mux_o_566;
wire mux_o_567;
wire mux_o_568;
wire mux_o_570;
wire mux_o_571;
wire mux_o_572;
wire mux_o_573;
wire mux_o_574;
wire mux_o_575;
wire mux_o_576;
wire mux_o_577;
wire mux_o_578;
wire mux_o_579;
wire mux_o_580;
wire mux_o_581;
wire mux_o_582;
wire mux_o_583;
wire mux_o_585;
wire mux_o_586;
wire mux_o_587;
wire mux_o_588;
wire mux_o_589;
wire mux_o_590;
wire mux_o_591;
wire mux_o_592;
wire mux_o_593;
wire mux_o_594;
wire mux_o_595;
wire mux_o_596;
wire mux_o_597;
wire mux_o_598;
wire mux_o_600;
wire mux_o_601;
wire mux_o_602;
wire mux_o_603;
wire mux_o_604;
wire mux_o_605;
wire mux_o_606;
wire mux_o_607;
wire mux_o_608;
wire mux_o_609;
wire mux_o_610;
wire mux_o_611;
wire mux_o_612;
wire mux_o_613;
wire mux_o_615;
wire mux_o_616;
wire mux_o_617;
wire mux_o_618;
wire mux_o_619;
wire mux_o_620;
wire mux_o_621;
wire mux_o_622;
wire mux_o_623;
wire mux_o_624;
wire mux_o_625;
wire mux_o_626;
wire mux_o_627;
wire mux_o_628;
wire mux_o_630;
wire mux_o_631;
wire mux_o_632;
wire mux_o_633;
wire mux_o_634;
wire mux_o_635;
wire mux_o_636;
wire mux_o_637;
wire mux_o_638;
wire mux_o_639;
wire mux_o_640;
wire mux_o_641;
wire mux_o_642;
wire mux_o_643;
wire mux_o_645;
wire mux_o_646;
wire mux_o_647;
wire mux_o_648;
wire mux_o_649;
wire mux_o_650;
wire mux_o_651;
wire mux_o_652;
wire mux_o_653;
wire mux_o_654;
wire mux_o_655;
wire mux_o_656;
wire mux_o_657;
wire mux_o_658;
wire mux_o_660;
wire mux_o_661;
wire mux_o_662;
wire mux_o_663;
wire mux_o_664;
wire mux_o_665;
wire mux_o_666;
wire mux_o_667;
wire mux_o_668;
wire mux_o_669;
wire mux_o_670;
wire mux_o_671;
wire mux_o_672;
wire mux_o_673;
wire mux_o_675;
wire mux_o_676;
wire mux_o_677;
wire mux_o_678;
wire mux_o_679;
wire mux_o_680;
wire mux_o_681;
wire mux_o_682;
wire mux_o_683;
wire mux_o_684;
wire mux_o_685;
wire mux_o_686;
wire mux_o_687;
wire mux_o_688;
wire mux_o_690;
wire mux_o_691;
wire mux_o_692;
wire mux_o_693;
wire mux_o_694;
wire mux_o_695;
wire mux_o_696;
wire mux_o_697;
wire mux_o_698;
wire mux_o_699;
wire mux_o_700;
wire mux_o_701;
wire mux_o_702;
wire mux_o_703;
wire mux_o_705;
wire mux_o_706;
wire mux_o_707;
wire mux_o_708;
wire mux_o_709;
wire mux_o_710;
wire mux_o_711;
wire mux_o_712;
wire mux_o_713;
wire mux_o_714;
wire mux_o_715;
wire mux_o_716;
wire mux_o_717;
wire mux_o_718;
wire mux_o_720;
wire mux_o_721;
wire mux_o_722;
wire mux_o_723;
wire mux_o_724;
wire mux_o_725;
wire mux_o_726;
wire mux_o_727;
wire mux_o_728;
wire mux_o_729;
wire mux_o_730;
wire mux_o_731;
wire mux_o_732;
wire mux_o_733;
wire mux_o_735;
wire mux_o_736;
wire mux_o_737;
wire mux_o_738;
wire mux_o_739;
wire mux_o_740;
wire mux_o_741;
wire mux_o_742;
wire mux_o_743;
wire mux_o_744;
wire mux_o_745;
wire mux_o_746;
wire mux_o_747;
wire mux_o_748;
wire mux_o_750;
wire mux_o_751;
wire mux_o_752;
wire mux_o_753;
wire mux_o_754;
wire mux_o_755;
wire mux_o_756;
wire mux_o_757;
wire mux_o_758;
wire mux_o_759;
wire mux_o_760;
wire mux_o_761;
wire mux_o_762;
wire mux_o_763;
wire mux_o_765;
wire mux_o_766;
wire mux_o_767;
wire mux_o_768;
wire mux_o_769;
wire mux_o_770;
wire mux_o_771;
wire mux_o_772;
wire mux_o_773;
wire mux_o_774;
wire mux_o_775;
wire mux_o_776;
wire mux_o_777;
wire mux_o_778;
wire mux_o_780;
wire mux_o_781;
wire mux_o_782;
wire mux_o_783;
wire mux_o_784;
wire mux_o_785;
wire mux_o_786;
wire mux_o_787;
wire mux_o_788;
wire mux_o_789;
wire mux_o_790;
wire mux_o_791;
wire mux_o_792;
wire mux_o_793;
wire mux_o_795;
wire mux_o_796;
wire mux_o_797;
wire mux_o_798;
wire mux_o_799;
wire mux_o_800;
wire mux_o_801;
wire mux_o_802;
wire mux_o_803;
wire mux_o_804;
wire mux_o_805;
wire mux_o_806;
wire mux_o_807;
wire mux_o_808;
wire mux_o_810;
wire mux_o_811;
wire mux_o_812;
wire mux_o_813;
wire mux_o_814;
wire mux_o_815;
wire mux_o_816;
wire mux_o_817;
wire mux_o_818;
wire mux_o_819;
wire mux_o_820;
wire mux_o_821;
wire mux_o_822;
wire mux_o_823;
wire mux_o_825;
wire mux_o_826;
wire mux_o_827;
wire mux_o_828;
wire mux_o_829;
wire mux_o_830;
wire mux_o_831;
wire mux_o_832;
wire mux_o_833;
wire mux_o_834;
wire mux_o_835;
wire mux_o_836;
wire mux_o_837;
wire mux_o_838;
wire mux_o_840;
wire mux_o_841;
wire mux_o_842;
wire mux_o_843;
wire mux_o_844;
wire mux_o_845;
wire mux_o_846;
wire mux_o_847;
wire mux_o_848;
wire mux_o_849;
wire mux_o_850;
wire mux_o_851;
wire mux_o_852;
wire mux_o_853;
wire mux_o_855;
wire mux_o_856;
wire mux_o_857;
wire mux_o_858;
wire mux_o_859;
wire mux_o_860;
wire mux_o_861;
wire mux_o_862;
wire mux_o_863;
wire mux_o_864;
wire mux_o_865;
wire mux_o_866;
wire mux_o_867;
wire mux_o_868;
wire mux_o_870;
wire mux_o_871;
wire mux_o_872;
wire mux_o_873;
wire mux_o_874;
wire mux_o_875;
wire mux_o_876;
wire mux_o_877;
wire mux_o_878;
wire mux_o_879;
wire mux_o_880;
wire mux_o_881;
wire mux_o_882;
wire mux_o_883;
wire mux_o_885;
wire mux_o_886;
wire mux_o_887;
wire mux_o_888;
wire mux_o_889;
wire mux_o_890;
wire mux_o_891;
wire mux_o_892;
wire mux_o_893;
wire mux_o_894;
wire mux_o_895;
wire mux_o_896;
wire mux_o_897;
wire mux_o_898;
wire mux_o_900;
wire mux_o_901;
wire mux_o_902;
wire mux_o_903;
wire mux_o_904;
wire mux_o_905;
wire mux_o_906;
wire mux_o_907;
wire mux_o_908;
wire mux_o_909;
wire mux_o_910;
wire mux_o_911;
wire mux_o_912;
wire mux_o_913;
wire mux_o_915;
wire mux_o_916;
wire mux_o_917;
wire mux_o_918;
wire mux_o_919;
wire mux_o_920;
wire mux_o_921;
wire mux_o_922;
wire mux_o_923;
wire mux_o_924;
wire mux_o_925;
wire mux_o_926;
wire mux_o_927;
wire mux_o_928;
wire mux_o_930;
wire mux_o_931;
wire mux_o_932;
wire mux_o_933;
wire mux_o_934;
wire mux_o_935;
wire mux_o_936;
wire mux_o_937;
wire mux_o_938;
wire mux_o_939;
wire mux_o_940;
wire mux_o_941;
wire mux_o_942;
wire mux_o_943;
wire mux_o_945;
wire mux_o_946;
wire mux_o_947;
wire mux_o_948;
wire mux_o_949;
wire mux_o_950;
wire mux_o_951;
wire mux_o_952;
wire mux_o_953;
wire mux_o_954;
wire mux_o_955;
wire mux_o_956;
wire mux_o_957;
wire mux_o_958;
wire cea_w;
wire ceb_w;
wire gw_gnd;

assign cea_w = ~wrea & cea;
assign ceb_w = ~wreb & ceb;
assign gw_gnd = 1'b0;

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13])
);
defparam lut_inst_0.INIT = 16'h0001;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13])
);
defparam lut_inst_1.INIT = 16'h0002;
LUT4 lut_inst_2 (
  .F(lut_f_2),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13])
);
defparam lut_inst_2.INIT = 16'h0004;
LUT4 lut_inst_3 (
  .F(lut_f_3),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13])
);
defparam lut_inst_3.INIT = 16'h0008;
LUT4 lut_inst_4 (
  .F(lut_f_4),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13])
);
defparam lut_inst_4.INIT = 16'h0010;
LUT4 lut_inst_5 (
  .F(lut_f_5),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13])
);
defparam lut_inst_5.INIT = 16'h0020;
LUT4 lut_inst_6 (
  .F(lut_f_6),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13])
);
defparam lut_inst_6.INIT = 16'h0040;
LUT4 lut_inst_7 (
  .F(lut_f_7),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13])
);
defparam lut_inst_7.INIT = 16'h0080;
LUT4 lut_inst_8 (
  .F(lut_f_8),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13])
);
defparam lut_inst_8.INIT = 16'h0100;
LUT4 lut_inst_9 (
  .F(lut_f_9),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13])
);
defparam lut_inst_9.INIT = 16'h0200;
LUT4 lut_inst_10 (
  .F(lut_f_10),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13])
);
defparam lut_inst_10.INIT = 16'h0400;
LUT4 lut_inst_11 (
  .F(lut_f_11),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13])
);
defparam lut_inst_11.INIT = 16'h0800;
LUT4 lut_inst_12 (
  .F(lut_f_12),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13])
);
defparam lut_inst_12.INIT = 16'h1000;
LUT4 lut_inst_13 (
  .F(lut_f_13),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13])
);
defparam lut_inst_13.INIT = 16'h2000;
LUT4 lut_inst_14 (
  .F(lut_f_14),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13])
);
defparam lut_inst_14.INIT = 16'h4000;
LUT4 lut_inst_15 (
  .F(lut_f_15),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13])
);
defparam lut_inst_15.INIT = 16'h8000;
LUT4 lut_inst_16 (
  .F(lut_f_16),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13])
);
defparam lut_inst_16.INIT = 16'h0001;
LUT4 lut_inst_17 (
  .F(lut_f_17),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13])
);
defparam lut_inst_17.INIT = 16'h0002;
LUT4 lut_inst_18 (
  .F(lut_f_18),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13])
);
defparam lut_inst_18.INIT = 16'h0004;
LUT4 lut_inst_19 (
  .F(lut_f_19),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13])
);
defparam lut_inst_19.INIT = 16'h0008;
LUT4 lut_inst_20 (
  .F(lut_f_20),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13])
);
defparam lut_inst_20.INIT = 16'h0010;
LUT4 lut_inst_21 (
  .F(lut_f_21),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13])
);
defparam lut_inst_21.INIT = 16'h0020;
LUT4 lut_inst_22 (
  .F(lut_f_22),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13])
);
defparam lut_inst_22.INIT = 16'h0040;
LUT4 lut_inst_23 (
  .F(lut_f_23),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13])
);
defparam lut_inst_23.INIT = 16'h0080;
LUT4 lut_inst_24 (
  .F(lut_f_24),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13])
);
defparam lut_inst_24.INIT = 16'h0100;
LUT4 lut_inst_25 (
  .F(lut_f_25),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13])
);
defparam lut_inst_25.INIT = 16'h0200;
LUT4 lut_inst_26 (
  .F(lut_f_26),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13])
);
defparam lut_inst_26.INIT = 16'h0400;
LUT4 lut_inst_27 (
  .F(lut_f_27),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13])
);
defparam lut_inst_27.INIT = 16'h0800;
LUT4 lut_inst_28 (
  .F(lut_f_28),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13])
);
defparam lut_inst_28.INIT = 16'h1000;
LUT4 lut_inst_29 (
  .F(lut_f_29),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13])
);
defparam lut_inst_29.INIT = 16'h2000;
LUT4 lut_inst_30 (
  .F(lut_f_30),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13])
);
defparam lut_inst_30.INIT = 16'h4000;
LUT4 lut_inst_31 (
  .F(lut_f_31),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13])
);
defparam lut_inst_31.INIT = 16'h8000;
DPB dpb_inst_0 (
    .DOA(dpb_inst_0_douta[15:0]),
    .DOB(dpb_inst_0_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_0}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_16}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_0.READ_MODE0 = 1'b0;
defparam dpb_inst_0.READ_MODE1 = 1'b0;
defparam dpb_inst_0.WRITE_MODE0 = 2'b00;
defparam dpb_inst_0.WRITE_MODE1 = 2'b00;
defparam dpb_inst_0.BIT_WIDTH_0 = 16;
defparam dpb_inst_0.BIT_WIDTH_1 = 16;
defparam dpb_inst_0.BLK_SEL_0 = 3'b001;
defparam dpb_inst_0.BLK_SEL_1 = 3'b001;
defparam dpb_inst_0.RESET_MODE = "SYNC";
defparam dpb_inst_0.INIT_RAM_00 = 256'h0000253B3B64323B5B1B0020253B3B64323B5B1B642564250078003C00040003;
defparam dpb_inst_0.INIT_RAM_01 = 256'h78666F6E006D303B323B5B1B006D303B323B5B1B96E20000253B3B64323B5B1B;
defparam dpb_inst_0.INIT_RAM_02 = 256'h544F73696E657275656D7475756F6667657475632073746E6572616520747475;
defparam dpb_inst_0.INIT_RAM_03 = 256'h000050432020732520206425250A0000313B38336D36353B5B1B000074616363;
defparam dpb_inst_0.INIT_RAM_04 = 256'h756F69776E697552325B5B1B313B38336D36353B5B1B3D534F54415200202020;
defparam dpb_inst_0.INIT_RAM_05 = 256'h444339383534313000002E29656D75736D20617263616F667475756F69687267;
defparam dpb_inst_0.INIT_RAM_06 = 256'h526052245224522452585324533853385258524C5324524C5258524C53380000;
defparam dpb_inst_0.INIT_RAM_07 = 256'h69D45A48595459545954598859585A48595859885A4859585958598859645964;
defparam dpb_inst_0.INIT_RAM_08 = 256'h6ECC6ECC6A7069EC69EC69EC6A686AD469D469D46A686A106AD46A106A686A10;
defparam dpb_inst_0.INIT_RAM_09 = 256'h0404030301006F546EC06EC06EC06EF06EC46F546EC46EF06F546EC46EC46EF0;
defparam dpb_inst_0.INIT_RAM_0A = 256'h0707070707070606060606060606060606060606060605050505050505050404;
defparam dpb_inst_0.INIT_RAM_0B = 256'h0808080808080707070707070707070707070707070707070707070707070707;
defparam dpb_inst_0.INIT_RAM_0C = 256'h0808080808080808080808080808080808080808080808080808080808080808;
defparam dpb_inst_0.INIT_RAM_0D = 256'h0000000000000808080808080808080808080808080808080808080808080808;
defparam dpb_inst_0.INIT_RAM_0E = 256'h000000000000126FCCCD000033330000CCCDCCCD999A0000000000000000F2CA;
defparam dpb_inst_0.INIT_RAM_0F = 256'h00000000000000000000666600000000000000000000000000000000CCCD999A;
defparam dpb_inst_0.INIT_RAM_10 = 256'h0000000079A743EC000000004000000000000000624DA9FC999A666600000000;
defparam dpb_inst_0.INIT_RAM_11 = 256'hAA3CC3A0384F38006DB7A3053255F1420000AA3BAAAB0000A570AA00CFDCC000;
defparam dpb_inst_0.INIT_RAM_12 = 256'h00004260F2CA0000000000000000AAAB0B61B355EA0EBB4CBE8C721872004260;
defparam dpb_inst_0.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_17 = 256'h001800480D1B7C017A0100000010000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_18 = 256'h0E44D844D644D444D244C8440270990A9707940592028108896C440005D43494;
defparam dpb_inst_0.INIT_RAM_19 = 256'h97079404810893038870440004F03A080018004C0D1B7C017A0100000010000B;
defparam dpb_inst_0.INIT_RAM_1A = 256'h000000000000000000000000000B0E44D944D744D544D344C944C10A030C990A;
defparam dpb_inst_0.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_1 (
    .DOA(dpb_inst_1_douta[15:0]),
    .DOB(dpb_inst_1_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_1}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_17}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_1.READ_MODE0 = 1'b0;
defparam dpb_inst_1.READ_MODE1 = 1'b0;
defparam dpb_inst_1.WRITE_MODE0 = 2'b00;
defparam dpb_inst_1.WRITE_MODE1 = 2'b00;
defparam dpb_inst_1.BIT_WIDTH_0 = 16;
defparam dpb_inst_1.BIT_WIDTH_1 = 16;
defparam dpb_inst_1.BLK_SEL_0 = 3'b001;
defparam dpb_inst_1.BLK_SEL_1 = 3'b001;
defparam dpb_inst_1.RESET_MODE = "SYNC";
defparam dpb_inst_1.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_2 (
    .DOA(dpb_inst_2_douta[15:0]),
    .DOB(dpb_inst_2_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_2}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_18}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_2.READ_MODE0 = 1'b0;
defparam dpb_inst_2.READ_MODE1 = 1'b0;
defparam dpb_inst_2.WRITE_MODE0 = 2'b00;
defparam dpb_inst_2.WRITE_MODE1 = 2'b00;
defparam dpb_inst_2.BIT_WIDTH_0 = 16;
defparam dpb_inst_2.BIT_WIDTH_1 = 16;
defparam dpb_inst_2.BLK_SEL_0 = 3'b001;
defparam dpb_inst_2.BLK_SEL_1 = 3'b001;
defparam dpb_inst_2.RESET_MODE = "SYNC";
defparam dpb_inst_2.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_3 (
    .DOA(dpb_inst_3_douta[15:0]),
    .DOB(dpb_inst_3_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_3}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_19}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_3.READ_MODE0 = 1'b0;
defparam dpb_inst_3.READ_MODE1 = 1'b0;
defparam dpb_inst_3.WRITE_MODE0 = 2'b00;
defparam dpb_inst_3.WRITE_MODE1 = 2'b00;
defparam dpb_inst_3.BIT_WIDTH_0 = 16;
defparam dpb_inst_3.BIT_WIDTH_1 = 16;
defparam dpb_inst_3.BLK_SEL_0 = 3'b001;
defparam dpb_inst_3.BLK_SEL_1 = 3'b001;
defparam dpb_inst_3.RESET_MODE = "SYNC";
defparam dpb_inst_3.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_4 (
    .DOA(dpb_inst_4_douta[15:0]),
    .DOB(dpb_inst_4_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_4}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_20}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_4.READ_MODE0 = 1'b0;
defparam dpb_inst_4.READ_MODE1 = 1'b0;
defparam dpb_inst_4.WRITE_MODE0 = 2'b00;
defparam dpb_inst_4.WRITE_MODE1 = 2'b00;
defparam dpb_inst_4.BIT_WIDTH_0 = 16;
defparam dpb_inst_4.BIT_WIDTH_1 = 16;
defparam dpb_inst_4.BLK_SEL_0 = 3'b001;
defparam dpb_inst_4.BLK_SEL_1 = 3'b001;
defparam dpb_inst_4.RESET_MODE = "SYNC";
defparam dpb_inst_4.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_5 (
    .DOA(dpb_inst_5_douta[15:0]),
    .DOB(dpb_inst_5_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_5}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_21}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_5.READ_MODE0 = 1'b0;
defparam dpb_inst_5.READ_MODE1 = 1'b0;
defparam dpb_inst_5.WRITE_MODE0 = 2'b00;
defparam dpb_inst_5.WRITE_MODE1 = 2'b00;
defparam dpb_inst_5.BIT_WIDTH_0 = 16;
defparam dpb_inst_5.BIT_WIDTH_1 = 16;
defparam dpb_inst_5.BLK_SEL_0 = 3'b001;
defparam dpb_inst_5.BLK_SEL_1 = 3'b001;
defparam dpb_inst_5.RESET_MODE = "SYNC";
defparam dpb_inst_5.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_5.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_6 (
    .DOA(dpb_inst_6_douta[15:0]),
    .DOB(dpb_inst_6_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_6}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_22}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_6.READ_MODE0 = 1'b0;
defparam dpb_inst_6.READ_MODE1 = 1'b0;
defparam dpb_inst_6.WRITE_MODE0 = 2'b00;
defparam dpb_inst_6.WRITE_MODE1 = 2'b00;
defparam dpb_inst_6.BIT_WIDTH_0 = 16;
defparam dpb_inst_6.BIT_WIDTH_1 = 16;
defparam dpb_inst_6.BLK_SEL_0 = 3'b001;
defparam dpb_inst_6.BLK_SEL_1 = 3'b001;
defparam dpb_inst_6.RESET_MODE = "SYNC";
defparam dpb_inst_6.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_6.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_7 (
    .DOA(dpb_inst_7_douta[15:0]),
    .DOB(dpb_inst_7_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_7}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_23}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_7.READ_MODE0 = 1'b0;
defparam dpb_inst_7.READ_MODE1 = 1'b0;
defparam dpb_inst_7.WRITE_MODE0 = 2'b00;
defparam dpb_inst_7.WRITE_MODE1 = 2'b00;
defparam dpb_inst_7.BIT_WIDTH_0 = 16;
defparam dpb_inst_7.BIT_WIDTH_1 = 16;
defparam dpb_inst_7.BLK_SEL_0 = 3'b001;
defparam dpb_inst_7.BLK_SEL_1 = 3'b001;
defparam dpb_inst_7.RESET_MODE = "SYNC";
defparam dpb_inst_7.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_7.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_8 (
    .DOA(dpb_inst_8_douta[15:0]),
    .DOB(dpb_inst_8_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_8}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_24}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_8.READ_MODE0 = 1'b0;
defparam dpb_inst_8.READ_MODE1 = 1'b0;
defparam dpb_inst_8.WRITE_MODE0 = 2'b00;
defparam dpb_inst_8.WRITE_MODE1 = 2'b00;
defparam dpb_inst_8.BIT_WIDTH_0 = 16;
defparam dpb_inst_8.BIT_WIDTH_1 = 16;
defparam dpb_inst_8.BLK_SEL_0 = 3'b001;
defparam dpb_inst_8.BLK_SEL_1 = 3'b001;
defparam dpb_inst_8.RESET_MODE = "SYNC";
defparam dpb_inst_8.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_8.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_9 (
    .DOA(dpb_inst_9_douta[15:0]),
    .DOB(dpb_inst_9_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_9}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_25}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_9.READ_MODE0 = 1'b0;
defparam dpb_inst_9.READ_MODE1 = 1'b0;
defparam dpb_inst_9.WRITE_MODE0 = 2'b00;
defparam dpb_inst_9.WRITE_MODE1 = 2'b00;
defparam dpb_inst_9.BIT_WIDTH_0 = 16;
defparam dpb_inst_9.BIT_WIDTH_1 = 16;
defparam dpb_inst_9.BLK_SEL_0 = 3'b001;
defparam dpb_inst_9.BLK_SEL_1 = 3'b001;
defparam dpb_inst_9.RESET_MODE = "SYNC";
defparam dpb_inst_9.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_10 (
    .DOA(dpb_inst_10_douta[15:0]),
    .DOB(dpb_inst_10_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_10}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_26}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_10.READ_MODE0 = 1'b0;
defparam dpb_inst_10.READ_MODE1 = 1'b0;
defparam dpb_inst_10.WRITE_MODE0 = 2'b00;
defparam dpb_inst_10.WRITE_MODE1 = 2'b00;
defparam dpb_inst_10.BIT_WIDTH_0 = 16;
defparam dpb_inst_10.BIT_WIDTH_1 = 16;
defparam dpb_inst_10.BLK_SEL_0 = 3'b001;
defparam dpb_inst_10.BLK_SEL_1 = 3'b001;
defparam dpb_inst_10.RESET_MODE = "SYNC";
defparam dpb_inst_10.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_10.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_11 (
    .DOA(dpb_inst_11_douta[15:0]),
    .DOB(dpb_inst_11_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_11}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_27}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_11.READ_MODE0 = 1'b0;
defparam dpb_inst_11.READ_MODE1 = 1'b0;
defparam dpb_inst_11.WRITE_MODE0 = 2'b00;
defparam dpb_inst_11.WRITE_MODE1 = 2'b00;
defparam dpb_inst_11.BIT_WIDTH_0 = 16;
defparam dpb_inst_11.BIT_WIDTH_1 = 16;
defparam dpb_inst_11.BLK_SEL_0 = 3'b001;
defparam dpb_inst_11.BLK_SEL_1 = 3'b001;
defparam dpb_inst_11.RESET_MODE = "SYNC";
defparam dpb_inst_11.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_11.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_12 (
    .DOA(dpb_inst_12_douta[15:0]),
    .DOB(dpb_inst_12_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_12}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_28}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_12.READ_MODE0 = 1'b0;
defparam dpb_inst_12.READ_MODE1 = 1'b0;
defparam dpb_inst_12.WRITE_MODE0 = 2'b00;
defparam dpb_inst_12.WRITE_MODE1 = 2'b00;
defparam dpb_inst_12.BIT_WIDTH_0 = 16;
defparam dpb_inst_12.BIT_WIDTH_1 = 16;
defparam dpb_inst_12.BLK_SEL_0 = 3'b001;
defparam dpb_inst_12.BLK_SEL_1 = 3'b001;
defparam dpb_inst_12.RESET_MODE = "SYNC";
defparam dpb_inst_12.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_12.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_13 (
    .DOA(dpb_inst_13_douta[15:0]),
    .DOB(dpb_inst_13_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_13}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_29}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_13.READ_MODE0 = 1'b0;
defparam dpb_inst_13.READ_MODE1 = 1'b0;
defparam dpb_inst_13.WRITE_MODE0 = 2'b00;
defparam dpb_inst_13.WRITE_MODE1 = 2'b00;
defparam dpb_inst_13.BIT_WIDTH_0 = 16;
defparam dpb_inst_13.BIT_WIDTH_1 = 16;
defparam dpb_inst_13.BLK_SEL_0 = 3'b001;
defparam dpb_inst_13.BLK_SEL_1 = 3'b001;
defparam dpb_inst_13.RESET_MODE = "SYNC";
defparam dpb_inst_13.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_13.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_14 (
    .DOA(dpb_inst_14_douta[15:0]),
    .DOB(dpb_inst_14_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_14}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_30}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_14.READ_MODE0 = 1'b0;
defparam dpb_inst_14.READ_MODE1 = 1'b0;
defparam dpb_inst_14.WRITE_MODE0 = 2'b00;
defparam dpb_inst_14.WRITE_MODE1 = 2'b00;
defparam dpb_inst_14.BIT_WIDTH_0 = 16;
defparam dpb_inst_14.BIT_WIDTH_1 = 16;
defparam dpb_inst_14.BLK_SEL_0 = 3'b001;
defparam dpb_inst_14.BLK_SEL_1 = 3'b001;
defparam dpb_inst_14.RESET_MODE = "SYNC";
defparam dpb_inst_14.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_14.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_15 (
    .DOA(dpb_inst_15_douta[15:0]),
    .DOB(dpb_inst_15_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_15}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_31}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_15.READ_MODE0 = 1'b0;
defparam dpb_inst_15.READ_MODE1 = 1'b0;
defparam dpb_inst_15.WRITE_MODE0 = 2'b00;
defparam dpb_inst_15.WRITE_MODE1 = 2'b00;
defparam dpb_inst_15.BIT_WIDTH_0 = 16;
defparam dpb_inst_15.BIT_WIDTH_1 = 16;
defparam dpb_inst_15.BLK_SEL_0 = 3'b001;
defparam dpb_inst_15.BLK_SEL_1 = 3'b001;
defparam dpb_inst_15.RESET_MODE = "SYNC";
defparam dpb_inst_15.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_15.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_16 (
    .DOA(dpb_inst_16_douta[31:16]),
    .DOB(dpb_inst_16_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_0}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_16}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_16.READ_MODE0 = 1'b0;
defparam dpb_inst_16.READ_MODE1 = 1'b0;
defparam dpb_inst_16.WRITE_MODE0 = 2'b00;
defparam dpb_inst_16.WRITE_MODE1 = 2'b00;
defparam dpb_inst_16.BIT_WIDTH_0 = 16;
defparam dpb_inst_16.BIT_WIDTH_1 = 16;
defparam dpb_inst_16.BLK_SEL_0 = 3'b001;
defparam dpb_inst_16.BLK_SEL_1 = 3'b001;
defparam dpb_inst_16.RESET_MODE = "SYNC";
defparam dpb_inst_16.INIT_RAM_00 = 256'h00006D646425253B383400006D646425253B38340000002E0000000000000000;
defparam dpb_inst_16.INIT_RAM_01 = 256'h6F2067200000303B303B38340000303B303B3833008300006D646425253B3833;
defparam dpb_inst_16.INIT_RAM_02 = 256'h61204E2020746D6573612820707420780029617263616920656D75736D287570;
defparam dpb_inst_16.INIT_RAM_03 = 256'h00003D490020202020202020786400006D35353B5B1B313B3834000029657275;
defparam dpb_inst_16.INIT_RAM_04 = 256'h2074687420676E6E004A1B486D35353B5B1B313B38340000454E535900002020;
defparam dpb_inst_16.INIT_RAM_05 = 256'h464542413736333200002E2E746E657261656574756320722820707420637061;
defparam dpb_inst_16.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
defparam dpb_inst_16.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_16.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_16.INIT_RAM_09 = 256'h040403030202FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_16.INIT_RAM_0A = 256'h0707070707070606060606060606060606060606060605050505050505050404;
defparam dpb_inst_16.INIT_RAM_0B = 256'h0808080808080707070707070707070707070707070707070707070707070707;
defparam dpb_inst_16.INIT_RAM_0C = 256'h0808080808080808080808080808080808080808080808080808080808080808;
defparam dpb_inst_16.INIT_RAM_0D = 256'hBF80437F3F800808080808080808080808080808080808080808080808080808;
defparam dpb_inst_16.INIT_RAM_0E = 256'h4000C180C0403A833F4C3F003F33447A3DCC3E4C3E99C1F0C120412040807149;
defparam dpb_inst_16.INIT_RAM_0F = 256'h41A0C1A0430E40A040E03F664040C190BF0042FA3FC0C140BFC042483ECC3F19;
defparam dpb_inst_16.INIT_RAM_10 = 256'h7F80FF803FF24FFE3FF00000408F00003FE000003F50D2F13FD93FE6C1C841F0;
defparam dpb_inst_16.INIT_RAM_11 = 256'h3338369D3F763F763EDB3E8B3E6C3E534B803FB83EAA3E8036EC3FB835D13F15;
defparam dpb_inst_16.INIT_RAM_12 = 256'h33008DA2F1494C00CB004B007FC03E2A3B36388A35DD333135BF3F313F310DA2;
defparam dpb_inst_16.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_17 = 256'h0000000000020101005200000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_18 = 256'h4400D944D744D544D344C944C10A030B98099506930488019603300E0000FFFF;
defparam dpb_inst_16.INIT_RAM_19 = 256'h98099506920196058902300E0000FFFF00000000000201010052000000000000;
defparam dpb_inst_16.INIT_RAM_1A = 256'h00000000000000000000000000004400DA44D844D644D444D244C84401209A0B;
defparam dpb_inst_16.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_16.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_17 (
    .DOA(dpb_inst_17_douta[31:16]),
    .DOB(dpb_inst_17_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_1}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_17}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_17.READ_MODE0 = 1'b0;
defparam dpb_inst_17.READ_MODE1 = 1'b0;
defparam dpb_inst_17.WRITE_MODE0 = 2'b00;
defparam dpb_inst_17.WRITE_MODE1 = 2'b00;
defparam dpb_inst_17.BIT_WIDTH_0 = 16;
defparam dpb_inst_17.BIT_WIDTH_1 = 16;
defparam dpb_inst_17.BLK_SEL_0 = 3'b001;
defparam dpb_inst_17.BLK_SEL_1 = 3'b001;
defparam dpb_inst_17.RESET_MODE = "SYNC";
defparam dpb_inst_17.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_17.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_18 (
    .DOA(dpb_inst_18_douta[31:16]),
    .DOB(dpb_inst_18_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_2}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_18}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_18.READ_MODE0 = 1'b0;
defparam dpb_inst_18.READ_MODE1 = 1'b0;
defparam dpb_inst_18.WRITE_MODE0 = 2'b00;
defparam dpb_inst_18.WRITE_MODE1 = 2'b00;
defparam dpb_inst_18.BIT_WIDTH_0 = 16;
defparam dpb_inst_18.BIT_WIDTH_1 = 16;
defparam dpb_inst_18.BLK_SEL_0 = 3'b001;
defparam dpb_inst_18.BLK_SEL_1 = 3'b001;
defparam dpb_inst_18.RESET_MODE = "SYNC";
defparam dpb_inst_18.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_18.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_19 (
    .DOA(dpb_inst_19_douta[31:16]),
    .DOB(dpb_inst_19_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_3}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_19}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_19.READ_MODE0 = 1'b0;
defparam dpb_inst_19.READ_MODE1 = 1'b0;
defparam dpb_inst_19.WRITE_MODE0 = 2'b00;
defparam dpb_inst_19.WRITE_MODE1 = 2'b00;
defparam dpb_inst_19.BIT_WIDTH_0 = 16;
defparam dpb_inst_19.BIT_WIDTH_1 = 16;
defparam dpb_inst_19.BLK_SEL_0 = 3'b001;
defparam dpb_inst_19.BLK_SEL_1 = 3'b001;
defparam dpb_inst_19.RESET_MODE = "SYNC";
defparam dpb_inst_19.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_19.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_20 (
    .DOA(dpb_inst_20_douta[31:16]),
    .DOB(dpb_inst_20_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_4}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_20}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_20.READ_MODE0 = 1'b0;
defparam dpb_inst_20.READ_MODE1 = 1'b0;
defparam dpb_inst_20.WRITE_MODE0 = 2'b00;
defparam dpb_inst_20.WRITE_MODE1 = 2'b00;
defparam dpb_inst_20.BIT_WIDTH_0 = 16;
defparam dpb_inst_20.BIT_WIDTH_1 = 16;
defparam dpb_inst_20.BLK_SEL_0 = 3'b001;
defparam dpb_inst_20.BLK_SEL_1 = 3'b001;
defparam dpb_inst_20.RESET_MODE = "SYNC";
defparam dpb_inst_20.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_20.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_21 (
    .DOA(dpb_inst_21_douta[31:16]),
    .DOB(dpb_inst_21_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_5}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_21}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_21.READ_MODE0 = 1'b0;
defparam dpb_inst_21.READ_MODE1 = 1'b0;
defparam dpb_inst_21.WRITE_MODE0 = 2'b00;
defparam dpb_inst_21.WRITE_MODE1 = 2'b00;
defparam dpb_inst_21.BIT_WIDTH_0 = 16;
defparam dpb_inst_21.BIT_WIDTH_1 = 16;
defparam dpb_inst_21.BLK_SEL_0 = 3'b001;
defparam dpb_inst_21.BLK_SEL_1 = 3'b001;
defparam dpb_inst_21.RESET_MODE = "SYNC";
defparam dpb_inst_21.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_21.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_22 (
    .DOA(dpb_inst_22_douta[31:16]),
    .DOB(dpb_inst_22_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_6}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_22}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_22.READ_MODE0 = 1'b0;
defparam dpb_inst_22.READ_MODE1 = 1'b0;
defparam dpb_inst_22.WRITE_MODE0 = 2'b00;
defparam dpb_inst_22.WRITE_MODE1 = 2'b00;
defparam dpb_inst_22.BIT_WIDTH_0 = 16;
defparam dpb_inst_22.BIT_WIDTH_1 = 16;
defparam dpb_inst_22.BLK_SEL_0 = 3'b001;
defparam dpb_inst_22.BLK_SEL_1 = 3'b001;
defparam dpb_inst_22.RESET_MODE = "SYNC";
defparam dpb_inst_22.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_22.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_23 (
    .DOA(dpb_inst_23_douta[31:16]),
    .DOB(dpb_inst_23_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_7}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_23}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_23.READ_MODE0 = 1'b0;
defparam dpb_inst_23.READ_MODE1 = 1'b0;
defparam dpb_inst_23.WRITE_MODE0 = 2'b00;
defparam dpb_inst_23.WRITE_MODE1 = 2'b00;
defparam dpb_inst_23.BIT_WIDTH_0 = 16;
defparam dpb_inst_23.BIT_WIDTH_1 = 16;
defparam dpb_inst_23.BLK_SEL_0 = 3'b001;
defparam dpb_inst_23.BLK_SEL_1 = 3'b001;
defparam dpb_inst_23.RESET_MODE = "SYNC";
defparam dpb_inst_23.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_23.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_24 (
    .DOA(dpb_inst_24_douta[31:16]),
    .DOB(dpb_inst_24_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_8}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_24}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_24.READ_MODE0 = 1'b0;
defparam dpb_inst_24.READ_MODE1 = 1'b0;
defparam dpb_inst_24.WRITE_MODE0 = 2'b00;
defparam dpb_inst_24.WRITE_MODE1 = 2'b00;
defparam dpb_inst_24.BIT_WIDTH_0 = 16;
defparam dpb_inst_24.BIT_WIDTH_1 = 16;
defparam dpb_inst_24.BLK_SEL_0 = 3'b001;
defparam dpb_inst_24.BLK_SEL_1 = 3'b001;
defparam dpb_inst_24.RESET_MODE = "SYNC";
defparam dpb_inst_24.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_25 (
    .DOA(dpb_inst_25_douta[31:16]),
    .DOB(dpb_inst_25_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_9}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_25}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_25.READ_MODE0 = 1'b0;
defparam dpb_inst_25.READ_MODE1 = 1'b0;
defparam dpb_inst_25.WRITE_MODE0 = 2'b00;
defparam dpb_inst_25.WRITE_MODE1 = 2'b00;
defparam dpb_inst_25.BIT_WIDTH_0 = 16;
defparam dpb_inst_25.BIT_WIDTH_1 = 16;
defparam dpb_inst_25.BLK_SEL_0 = 3'b001;
defparam dpb_inst_25.BLK_SEL_1 = 3'b001;
defparam dpb_inst_25.RESET_MODE = "SYNC";
defparam dpb_inst_25.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_26 (
    .DOA(dpb_inst_26_douta[31:16]),
    .DOB(dpb_inst_26_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_10}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_26}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_26.READ_MODE0 = 1'b0;
defparam dpb_inst_26.READ_MODE1 = 1'b0;
defparam dpb_inst_26.WRITE_MODE0 = 2'b00;
defparam dpb_inst_26.WRITE_MODE1 = 2'b00;
defparam dpb_inst_26.BIT_WIDTH_0 = 16;
defparam dpb_inst_26.BIT_WIDTH_1 = 16;
defparam dpb_inst_26.BLK_SEL_0 = 3'b001;
defparam dpb_inst_26.BLK_SEL_1 = 3'b001;
defparam dpb_inst_26.RESET_MODE = "SYNC";
defparam dpb_inst_26.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_27 (
    .DOA(dpb_inst_27_douta[31:16]),
    .DOB(dpb_inst_27_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_11}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_27}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_27.READ_MODE0 = 1'b0;
defparam dpb_inst_27.READ_MODE1 = 1'b0;
defparam dpb_inst_27.WRITE_MODE0 = 2'b00;
defparam dpb_inst_27.WRITE_MODE1 = 2'b00;
defparam dpb_inst_27.BIT_WIDTH_0 = 16;
defparam dpb_inst_27.BIT_WIDTH_1 = 16;
defparam dpb_inst_27.BLK_SEL_0 = 3'b001;
defparam dpb_inst_27.BLK_SEL_1 = 3'b001;
defparam dpb_inst_27.RESET_MODE = "SYNC";
defparam dpb_inst_27.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_28 (
    .DOA(dpb_inst_28_douta[31:16]),
    .DOB(dpb_inst_28_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_12}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_28}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_28.READ_MODE0 = 1'b0;
defparam dpb_inst_28.READ_MODE1 = 1'b0;
defparam dpb_inst_28.WRITE_MODE0 = 2'b00;
defparam dpb_inst_28.WRITE_MODE1 = 2'b00;
defparam dpb_inst_28.BIT_WIDTH_0 = 16;
defparam dpb_inst_28.BIT_WIDTH_1 = 16;
defparam dpb_inst_28.BLK_SEL_0 = 3'b001;
defparam dpb_inst_28.BLK_SEL_1 = 3'b001;
defparam dpb_inst_28.RESET_MODE = "SYNC";
defparam dpb_inst_28.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_29 (
    .DOA(dpb_inst_29_douta[31:16]),
    .DOB(dpb_inst_29_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_13}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_29}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_29.READ_MODE0 = 1'b0;
defparam dpb_inst_29.READ_MODE1 = 1'b0;
defparam dpb_inst_29.WRITE_MODE0 = 2'b00;
defparam dpb_inst_29.WRITE_MODE1 = 2'b00;
defparam dpb_inst_29.BIT_WIDTH_0 = 16;
defparam dpb_inst_29.BIT_WIDTH_1 = 16;
defparam dpb_inst_29.BLK_SEL_0 = 3'b001;
defparam dpb_inst_29.BLK_SEL_1 = 3'b001;
defparam dpb_inst_29.RESET_MODE = "SYNC";
defparam dpb_inst_29.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_29.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_30 (
    .DOA(dpb_inst_30_douta[31:16]),
    .DOB(dpb_inst_30_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_14}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_30}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_30.READ_MODE0 = 1'b0;
defparam dpb_inst_30.READ_MODE1 = 1'b0;
defparam dpb_inst_30.WRITE_MODE0 = 2'b00;
defparam dpb_inst_30.WRITE_MODE1 = 2'b00;
defparam dpb_inst_30.BIT_WIDTH_0 = 16;
defparam dpb_inst_30.BIT_WIDTH_1 = 16;
defparam dpb_inst_30.BLK_SEL_0 = 3'b001;
defparam dpb_inst_30.BLK_SEL_1 = 3'b001;
defparam dpb_inst_30.RESET_MODE = "SYNC";
defparam dpb_inst_30.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_30.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_31 (
    .DOA(dpb_inst_31_douta[31:16]),
    .DOB(dpb_inst_31_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_15}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_31}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_31.READ_MODE0 = 1'b0;
defparam dpb_inst_31.READ_MODE1 = 1'b0;
defparam dpb_inst_31.WRITE_MODE0 = 2'b00;
defparam dpb_inst_31.WRITE_MODE1 = 2'b00;
defparam dpb_inst_31.BIT_WIDTH_0 = 16;
defparam dpb_inst_31.BIT_WIDTH_1 = 16;
defparam dpb_inst_31.BLK_SEL_0 = 3'b001;
defparam dpb_inst_31.BLK_SEL_1 = 3'b001;
defparam dpb_inst_31.RESET_MODE = "SYNC";
defparam dpb_inst_31.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_31.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DFFRE dff_inst_0 (
  .Q(dff_q_0),
  .D(ada[13]),
  .CLK(clka),
  .CE(cea_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_1 (
  .Q(dff_q_1),
  .D(ada[12]),
  .CLK(clka),
  .CE(cea_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_2 (
  .Q(dff_q_2),
  .D(ada[11]),
  .CLK(clka),
  .CE(cea_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_3 (
  .Q(dff_q_3),
  .D(ada[10]),
  .CLK(clka),
  .CE(cea_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_4 (
  .Q(dff_q_4),
  .D(adb[13]),
  .CLK(clkb),
  .CE(ceb_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_5 (
  .Q(dff_q_5),
  .D(adb[12]),
  .CLK(clkb),
  .CE(ceb_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_6 (
  .Q(dff_q_6),
  .D(adb[11]),
  .CLK(clkb),
  .CE(ceb_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_7 (
  .Q(dff_q_7),
  .D(adb[10]),
  .CLK(clkb),
  .CE(ceb_w),
  .RESET(gw_gnd)
);
MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(dpb_inst_0_douta[0]),
  .I1(dpb_inst_1_douta[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(dpb_inst_2_douta[0]),
  .I1(dpb_inst_3_douta[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(dpb_inst_4_douta[0]),
  .I1(dpb_inst_5_douta[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(dpb_inst_6_douta[0]),
  .I1(dpb_inst_7_douta[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(dpb_inst_8_douta[0]),
  .I1(dpb_inst_9_douta[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(dpb_inst_10_douta[0]),
  .I1(dpb_inst_11_douta[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(dpb_inst_12_douta[0]),
  .I1(dpb_inst_13_douta[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_7 (
  .O(mux_o_7),
  .I0(dpb_inst_14_douta[0]),
  .I1(dpb_inst_15_douta[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(dff_q_2)
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(dff_q_2)
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(dff_q_2)
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(mux_o_6),
  .I1(mux_o_7),
  .S0(dff_q_2)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(mux_o_8),
  .I1(mux_o_9),
  .S0(dff_q_1)
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(mux_o_10),
  .I1(mux_o_11),
  .S0(dff_q_1)
);
MUX2 mux_inst_14 (
  .O(douta[0]),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(dff_q_0)
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(dpb_inst_0_douta[1]),
  .I1(dpb_inst_1_douta[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(dpb_inst_2_douta[1]),
  .I1(dpb_inst_3_douta[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(dpb_inst_4_douta[1]),
  .I1(dpb_inst_5_douta[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(dpb_inst_6_douta[1]),
  .I1(dpb_inst_7_douta[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_19 (
  .O(mux_o_19),
  .I0(dpb_inst_8_douta[1]),
  .I1(dpb_inst_9_douta[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_20 (
  .O(mux_o_20),
  .I0(dpb_inst_10_douta[1]),
  .I1(dpb_inst_11_douta[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(dpb_inst_12_douta[1]),
  .I1(dpb_inst_13_douta[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_22 (
  .O(mux_o_22),
  .I0(dpb_inst_14_douta[1]),
  .I1(dpb_inst_15_douta[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_23 (
  .O(mux_o_23),
  .I0(mux_o_15),
  .I1(mux_o_16),
  .S0(dff_q_2)
);
MUX2 mux_inst_24 (
  .O(mux_o_24),
  .I0(mux_o_17),
  .I1(mux_o_18),
  .S0(dff_q_2)
);
MUX2 mux_inst_25 (
  .O(mux_o_25),
  .I0(mux_o_19),
  .I1(mux_o_20),
  .S0(dff_q_2)
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(mux_o_21),
  .I1(mux_o_22),
  .S0(dff_q_2)
);
MUX2 mux_inst_27 (
  .O(mux_o_27),
  .I0(mux_o_23),
  .I1(mux_o_24),
  .S0(dff_q_1)
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(mux_o_25),
  .I1(mux_o_26),
  .S0(dff_q_1)
);
MUX2 mux_inst_29 (
  .O(douta[1]),
  .I0(mux_o_27),
  .I1(mux_o_28),
  .S0(dff_q_0)
);
MUX2 mux_inst_30 (
  .O(mux_o_30),
  .I0(dpb_inst_0_douta[2]),
  .I1(dpb_inst_1_douta[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(dpb_inst_2_douta[2]),
  .I1(dpb_inst_3_douta[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(dpb_inst_4_douta[2]),
  .I1(dpb_inst_5_douta[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(dpb_inst_6_douta[2]),
  .I1(dpb_inst_7_douta[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(dpb_inst_8_douta[2]),
  .I1(dpb_inst_9_douta[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(dpb_inst_10_douta[2]),
  .I1(dpb_inst_11_douta[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(dpb_inst_12_douta[2]),
  .I1(dpb_inst_13_douta[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_37 (
  .O(mux_o_37),
  .I0(dpb_inst_14_douta[2]),
  .I1(dpb_inst_15_douta[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_38 (
  .O(mux_o_38),
  .I0(mux_o_30),
  .I1(mux_o_31),
  .S0(dff_q_2)
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(mux_o_32),
  .I1(mux_o_33),
  .S0(dff_q_2)
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(mux_o_34),
  .I1(mux_o_35),
  .S0(dff_q_2)
);
MUX2 mux_inst_41 (
  .O(mux_o_41),
  .I0(mux_o_36),
  .I1(mux_o_37),
  .S0(dff_q_2)
);
MUX2 mux_inst_42 (
  .O(mux_o_42),
  .I0(mux_o_38),
  .I1(mux_o_39),
  .S0(dff_q_1)
);
MUX2 mux_inst_43 (
  .O(mux_o_43),
  .I0(mux_o_40),
  .I1(mux_o_41),
  .S0(dff_q_1)
);
MUX2 mux_inst_44 (
  .O(douta[2]),
  .I0(mux_o_42),
  .I1(mux_o_43),
  .S0(dff_q_0)
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(dpb_inst_0_douta[3]),
  .I1(dpb_inst_1_douta[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(dpb_inst_2_douta[3]),
  .I1(dpb_inst_3_douta[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_47 (
  .O(mux_o_47),
  .I0(dpb_inst_4_douta[3]),
  .I1(dpb_inst_5_douta[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_48 (
  .O(mux_o_48),
  .I0(dpb_inst_6_douta[3]),
  .I1(dpb_inst_7_douta[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_49 (
  .O(mux_o_49),
  .I0(dpb_inst_8_douta[3]),
  .I1(dpb_inst_9_douta[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(dpb_inst_10_douta[3]),
  .I1(dpb_inst_11_douta[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_51 (
  .O(mux_o_51),
  .I0(dpb_inst_12_douta[3]),
  .I1(dpb_inst_13_douta[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_52 (
  .O(mux_o_52),
  .I0(dpb_inst_14_douta[3]),
  .I1(dpb_inst_15_douta[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_53 (
  .O(mux_o_53),
  .I0(mux_o_45),
  .I1(mux_o_46),
  .S0(dff_q_2)
);
MUX2 mux_inst_54 (
  .O(mux_o_54),
  .I0(mux_o_47),
  .I1(mux_o_48),
  .S0(dff_q_2)
);
MUX2 mux_inst_55 (
  .O(mux_o_55),
  .I0(mux_o_49),
  .I1(mux_o_50),
  .S0(dff_q_2)
);
MUX2 mux_inst_56 (
  .O(mux_o_56),
  .I0(mux_o_51),
  .I1(mux_o_52),
  .S0(dff_q_2)
);
MUX2 mux_inst_57 (
  .O(mux_o_57),
  .I0(mux_o_53),
  .I1(mux_o_54),
  .S0(dff_q_1)
);
MUX2 mux_inst_58 (
  .O(mux_o_58),
  .I0(mux_o_55),
  .I1(mux_o_56),
  .S0(dff_q_1)
);
MUX2 mux_inst_59 (
  .O(douta[3]),
  .I0(mux_o_57),
  .I1(mux_o_58),
  .S0(dff_q_0)
);
MUX2 mux_inst_60 (
  .O(mux_o_60),
  .I0(dpb_inst_0_douta[4]),
  .I1(dpb_inst_1_douta[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_61 (
  .O(mux_o_61),
  .I0(dpb_inst_2_douta[4]),
  .I1(dpb_inst_3_douta[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_62 (
  .O(mux_o_62),
  .I0(dpb_inst_4_douta[4]),
  .I1(dpb_inst_5_douta[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_63 (
  .O(mux_o_63),
  .I0(dpb_inst_6_douta[4]),
  .I1(dpb_inst_7_douta[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_64 (
  .O(mux_o_64),
  .I0(dpb_inst_8_douta[4]),
  .I1(dpb_inst_9_douta[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_65 (
  .O(mux_o_65),
  .I0(dpb_inst_10_douta[4]),
  .I1(dpb_inst_11_douta[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_66 (
  .O(mux_o_66),
  .I0(dpb_inst_12_douta[4]),
  .I1(dpb_inst_13_douta[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_67 (
  .O(mux_o_67),
  .I0(dpb_inst_14_douta[4]),
  .I1(dpb_inst_15_douta[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_68 (
  .O(mux_o_68),
  .I0(mux_o_60),
  .I1(mux_o_61),
  .S0(dff_q_2)
);
MUX2 mux_inst_69 (
  .O(mux_o_69),
  .I0(mux_o_62),
  .I1(mux_o_63),
  .S0(dff_q_2)
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(mux_o_64),
  .I1(mux_o_65),
  .S0(dff_q_2)
);
MUX2 mux_inst_71 (
  .O(mux_o_71),
  .I0(mux_o_66),
  .I1(mux_o_67),
  .S0(dff_q_2)
);
MUX2 mux_inst_72 (
  .O(mux_o_72),
  .I0(mux_o_68),
  .I1(mux_o_69),
  .S0(dff_q_1)
);
MUX2 mux_inst_73 (
  .O(mux_o_73),
  .I0(mux_o_70),
  .I1(mux_o_71),
  .S0(dff_q_1)
);
MUX2 mux_inst_74 (
  .O(douta[4]),
  .I0(mux_o_72),
  .I1(mux_o_73),
  .S0(dff_q_0)
);
MUX2 mux_inst_75 (
  .O(mux_o_75),
  .I0(dpb_inst_0_douta[5]),
  .I1(dpb_inst_1_douta[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_76 (
  .O(mux_o_76),
  .I0(dpb_inst_2_douta[5]),
  .I1(dpb_inst_3_douta[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_77 (
  .O(mux_o_77),
  .I0(dpb_inst_4_douta[5]),
  .I1(dpb_inst_5_douta[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(dpb_inst_6_douta[5]),
  .I1(dpb_inst_7_douta[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(dpb_inst_8_douta[5]),
  .I1(dpb_inst_9_douta[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_80 (
  .O(mux_o_80),
  .I0(dpb_inst_10_douta[5]),
  .I1(dpb_inst_11_douta[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_81 (
  .O(mux_o_81),
  .I0(dpb_inst_12_douta[5]),
  .I1(dpb_inst_13_douta[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(dpb_inst_14_douta[5]),
  .I1(dpb_inst_15_douta[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_83 (
  .O(mux_o_83),
  .I0(mux_o_75),
  .I1(mux_o_76),
  .S0(dff_q_2)
);
MUX2 mux_inst_84 (
  .O(mux_o_84),
  .I0(mux_o_77),
  .I1(mux_o_78),
  .S0(dff_q_2)
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(mux_o_79),
  .I1(mux_o_80),
  .S0(dff_q_2)
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(mux_o_81),
  .I1(mux_o_82),
  .S0(dff_q_2)
);
MUX2 mux_inst_87 (
  .O(mux_o_87),
  .I0(mux_o_83),
  .I1(mux_o_84),
  .S0(dff_q_1)
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(mux_o_85),
  .I1(mux_o_86),
  .S0(dff_q_1)
);
MUX2 mux_inst_89 (
  .O(douta[5]),
  .I0(mux_o_87),
  .I1(mux_o_88),
  .S0(dff_q_0)
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(dpb_inst_0_douta[6]),
  .I1(dpb_inst_1_douta[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(dpb_inst_2_douta[6]),
  .I1(dpb_inst_3_douta[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_92 (
  .O(mux_o_92),
  .I0(dpb_inst_4_douta[6]),
  .I1(dpb_inst_5_douta[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(dpb_inst_6_douta[6]),
  .I1(dpb_inst_7_douta[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_94 (
  .O(mux_o_94),
  .I0(dpb_inst_8_douta[6]),
  .I1(dpb_inst_9_douta[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_95 (
  .O(mux_o_95),
  .I0(dpb_inst_10_douta[6]),
  .I1(dpb_inst_11_douta[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_96 (
  .O(mux_o_96),
  .I0(dpb_inst_12_douta[6]),
  .I1(dpb_inst_13_douta[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_97 (
  .O(mux_o_97),
  .I0(dpb_inst_14_douta[6]),
  .I1(dpb_inst_15_douta[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_98 (
  .O(mux_o_98),
  .I0(mux_o_90),
  .I1(mux_o_91),
  .S0(dff_q_2)
);
MUX2 mux_inst_99 (
  .O(mux_o_99),
  .I0(mux_o_92),
  .I1(mux_o_93),
  .S0(dff_q_2)
);
MUX2 mux_inst_100 (
  .O(mux_o_100),
  .I0(mux_o_94),
  .I1(mux_o_95),
  .S0(dff_q_2)
);
MUX2 mux_inst_101 (
  .O(mux_o_101),
  .I0(mux_o_96),
  .I1(mux_o_97),
  .S0(dff_q_2)
);
MUX2 mux_inst_102 (
  .O(mux_o_102),
  .I0(mux_o_98),
  .I1(mux_o_99),
  .S0(dff_q_1)
);
MUX2 mux_inst_103 (
  .O(mux_o_103),
  .I0(mux_o_100),
  .I1(mux_o_101),
  .S0(dff_q_1)
);
MUX2 mux_inst_104 (
  .O(douta[6]),
  .I0(mux_o_102),
  .I1(mux_o_103),
  .S0(dff_q_0)
);
MUX2 mux_inst_105 (
  .O(mux_o_105),
  .I0(dpb_inst_0_douta[7]),
  .I1(dpb_inst_1_douta[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_106 (
  .O(mux_o_106),
  .I0(dpb_inst_2_douta[7]),
  .I1(dpb_inst_3_douta[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(dpb_inst_4_douta[7]),
  .I1(dpb_inst_5_douta[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(dpb_inst_6_douta[7]),
  .I1(dpb_inst_7_douta[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(dpb_inst_8_douta[7]),
  .I1(dpb_inst_9_douta[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_110 (
  .O(mux_o_110),
  .I0(dpb_inst_10_douta[7]),
  .I1(dpb_inst_11_douta[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_111 (
  .O(mux_o_111),
  .I0(dpb_inst_12_douta[7]),
  .I1(dpb_inst_13_douta[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(dpb_inst_14_douta[7]),
  .I1(dpb_inst_15_douta[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_113 (
  .O(mux_o_113),
  .I0(mux_o_105),
  .I1(mux_o_106),
  .S0(dff_q_2)
);
MUX2 mux_inst_114 (
  .O(mux_o_114),
  .I0(mux_o_107),
  .I1(mux_o_108),
  .S0(dff_q_2)
);
MUX2 mux_inst_115 (
  .O(mux_o_115),
  .I0(mux_o_109),
  .I1(mux_o_110),
  .S0(dff_q_2)
);
MUX2 mux_inst_116 (
  .O(mux_o_116),
  .I0(mux_o_111),
  .I1(mux_o_112),
  .S0(dff_q_2)
);
MUX2 mux_inst_117 (
  .O(mux_o_117),
  .I0(mux_o_113),
  .I1(mux_o_114),
  .S0(dff_q_1)
);
MUX2 mux_inst_118 (
  .O(mux_o_118),
  .I0(mux_o_115),
  .I1(mux_o_116),
  .S0(dff_q_1)
);
MUX2 mux_inst_119 (
  .O(douta[7]),
  .I0(mux_o_117),
  .I1(mux_o_118),
  .S0(dff_q_0)
);
MUX2 mux_inst_120 (
  .O(mux_o_120),
  .I0(dpb_inst_0_douta[8]),
  .I1(dpb_inst_1_douta[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_121 (
  .O(mux_o_121),
  .I0(dpb_inst_2_douta[8]),
  .I1(dpb_inst_3_douta[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_122 (
  .O(mux_o_122),
  .I0(dpb_inst_4_douta[8]),
  .I1(dpb_inst_5_douta[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_123 (
  .O(mux_o_123),
  .I0(dpb_inst_6_douta[8]),
  .I1(dpb_inst_7_douta[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_124 (
  .O(mux_o_124),
  .I0(dpb_inst_8_douta[8]),
  .I1(dpb_inst_9_douta[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_125 (
  .O(mux_o_125),
  .I0(dpb_inst_10_douta[8]),
  .I1(dpb_inst_11_douta[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_126 (
  .O(mux_o_126),
  .I0(dpb_inst_12_douta[8]),
  .I1(dpb_inst_13_douta[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_127 (
  .O(mux_o_127),
  .I0(dpb_inst_14_douta[8]),
  .I1(dpb_inst_15_douta[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_128 (
  .O(mux_o_128),
  .I0(mux_o_120),
  .I1(mux_o_121),
  .S0(dff_q_2)
);
MUX2 mux_inst_129 (
  .O(mux_o_129),
  .I0(mux_o_122),
  .I1(mux_o_123),
  .S0(dff_q_2)
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(mux_o_124),
  .I1(mux_o_125),
  .S0(dff_q_2)
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(mux_o_126),
  .I1(mux_o_127),
  .S0(dff_q_2)
);
MUX2 mux_inst_132 (
  .O(mux_o_132),
  .I0(mux_o_128),
  .I1(mux_o_129),
  .S0(dff_q_1)
);
MUX2 mux_inst_133 (
  .O(mux_o_133),
  .I0(mux_o_130),
  .I1(mux_o_131),
  .S0(dff_q_1)
);
MUX2 mux_inst_134 (
  .O(douta[8]),
  .I0(mux_o_132),
  .I1(mux_o_133),
  .S0(dff_q_0)
);
MUX2 mux_inst_135 (
  .O(mux_o_135),
  .I0(dpb_inst_0_douta[9]),
  .I1(dpb_inst_1_douta[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_136 (
  .O(mux_o_136),
  .I0(dpb_inst_2_douta[9]),
  .I1(dpb_inst_3_douta[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_137 (
  .O(mux_o_137),
  .I0(dpb_inst_4_douta[9]),
  .I1(dpb_inst_5_douta[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_138 (
  .O(mux_o_138),
  .I0(dpb_inst_6_douta[9]),
  .I1(dpb_inst_7_douta[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_139 (
  .O(mux_o_139),
  .I0(dpb_inst_8_douta[9]),
  .I1(dpb_inst_9_douta[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_140 (
  .O(mux_o_140),
  .I0(dpb_inst_10_douta[9]),
  .I1(dpb_inst_11_douta[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_141 (
  .O(mux_o_141),
  .I0(dpb_inst_12_douta[9]),
  .I1(dpb_inst_13_douta[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_142 (
  .O(mux_o_142),
  .I0(dpb_inst_14_douta[9]),
  .I1(dpb_inst_15_douta[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_143 (
  .O(mux_o_143),
  .I0(mux_o_135),
  .I1(mux_o_136),
  .S0(dff_q_2)
);
MUX2 mux_inst_144 (
  .O(mux_o_144),
  .I0(mux_o_137),
  .I1(mux_o_138),
  .S0(dff_q_2)
);
MUX2 mux_inst_145 (
  .O(mux_o_145),
  .I0(mux_o_139),
  .I1(mux_o_140),
  .S0(dff_q_2)
);
MUX2 mux_inst_146 (
  .O(mux_o_146),
  .I0(mux_o_141),
  .I1(mux_o_142),
  .S0(dff_q_2)
);
MUX2 mux_inst_147 (
  .O(mux_o_147),
  .I0(mux_o_143),
  .I1(mux_o_144),
  .S0(dff_q_1)
);
MUX2 mux_inst_148 (
  .O(mux_o_148),
  .I0(mux_o_145),
  .I1(mux_o_146),
  .S0(dff_q_1)
);
MUX2 mux_inst_149 (
  .O(douta[9]),
  .I0(mux_o_147),
  .I1(mux_o_148),
  .S0(dff_q_0)
);
MUX2 mux_inst_150 (
  .O(mux_o_150),
  .I0(dpb_inst_0_douta[10]),
  .I1(dpb_inst_1_douta[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_151 (
  .O(mux_o_151),
  .I0(dpb_inst_2_douta[10]),
  .I1(dpb_inst_3_douta[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_152 (
  .O(mux_o_152),
  .I0(dpb_inst_4_douta[10]),
  .I1(dpb_inst_5_douta[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_153 (
  .O(mux_o_153),
  .I0(dpb_inst_6_douta[10]),
  .I1(dpb_inst_7_douta[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_154 (
  .O(mux_o_154),
  .I0(dpb_inst_8_douta[10]),
  .I1(dpb_inst_9_douta[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_155 (
  .O(mux_o_155),
  .I0(dpb_inst_10_douta[10]),
  .I1(dpb_inst_11_douta[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_156 (
  .O(mux_o_156),
  .I0(dpb_inst_12_douta[10]),
  .I1(dpb_inst_13_douta[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_157 (
  .O(mux_o_157),
  .I0(dpb_inst_14_douta[10]),
  .I1(dpb_inst_15_douta[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_158 (
  .O(mux_o_158),
  .I0(mux_o_150),
  .I1(mux_o_151),
  .S0(dff_q_2)
);
MUX2 mux_inst_159 (
  .O(mux_o_159),
  .I0(mux_o_152),
  .I1(mux_o_153),
  .S0(dff_q_2)
);
MUX2 mux_inst_160 (
  .O(mux_o_160),
  .I0(mux_o_154),
  .I1(mux_o_155),
  .S0(dff_q_2)
);
MUX2 mux_inst_161 (
  .O(mux_o_161),
  .I0(mux_o_156),
  .I1(mux_o_157),
  .S0(dff_q_2)
);
MUX2 mux_inst_162 (
  .O(mux_o_162),
  .I0(mux_o_158),
  .I1(mux_o_159),
  .S0(dff_q_1)
);
MUX2 mux_inst_163 (
  .O(mux_o_163),
  .I0(mux_o_160),
  .I1(mux_o_161),
  .S0(dff_q_1)
);
MUX2 mux_inst_164 (
  .O(douta[10]),
  .I0(mux_o_162),
  .I1(mux_o_163),
  .S0(dff_q_0)
);
MUX2 mux_inst_165 (
  .O(mux_o_165),
  .I0(dpb_inst_0_douta[11]),
  .I1(dpb_inst_1_douta[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_166 (
  .O(mux_o_166),
  .I0(dpb_inst_2_douta[11]),
  .I1(dpb_inst_3_douta[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_167 (
  .O(mux_o_167),
  .I0(dpb_inst_4_douta[11]),
  .I1(dpb_inst_5_douta[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_168 (
  .O(mux_o_168),
  .I0(dpb_inst_6_douta[11]),
  .I1(dpb_inst_7_douta[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_169 (
  .O(mux_o_169),
  .I0(dpb_inst_8_douta[11]),
  .I1(dpb_inst_9_douta[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_170 (
  .O(mux_o_170),
  .I0(dpb_inst_10_douta[11]),
  .I1(dpb_inst_11_douta[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_171 (
  .O(mux_o_171),
  .I0(dpb_inst_12_douta[11]),
  .I1(dpb_inst_13_douta[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_172 (
  .O(mux_o_172),
  .I0(dpb_inst_14_douta[11]),
  .I1(dpb_inst_15_douta[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_173 (
  .O(mux_o_173),
  .I0(mux_o_165),
  .I1(mux_o_166),
  .S0(dff_q_2)
);
MUX2 mux_inst_174 (
  .O(mux_o_174),
  .I0(mux_o_167),
  .I1(mux_o_168),
  .S0(dff_q_2)
);
MUX2 mux_inst_175 (
  .O(mux_o_175),
  .I0(mux_o_169),
  .I1(mux_o_170),
  .S0(dff_q_2)
);
MUX2 mux_inst_176 (
  .O(mux_o_176),
  .I0(mux_o_171),
  .I1(mux_o_172),
  .S0(dff_q_2)
);
MUX2 mux_inst_177 (
  .O(mux_o_177),
  .I0(mux_o_173),
  .I1(mux_o_174),
  .S0(dff_q_1)
);
MUX2 mux_inst_178 (
  .O(mux_o_178),
  .I0(mux_o_175),
  .I1(mux_o_176),
  .S0(dff_q_1)
);
MUX2 mux_inst_179 (
  .O(douta[11]),
  .I0(mux_o_177),
  .I1(mux_o_178),
  .S0(dff_q_0)
);
MUX2 mux_inst_180 (
  .O(mux_o_180),
  .I0(dpb_inst_0_douta[12]),
  .I1(dpb_inst_1_douta[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_181 (
  .O(mux_o_181),
  .I0(dpb_inst_2_douta[12]),
  .I1(dpb_inst_3_douta[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(dpb_inst_4_douta[12]),
  .I1(dpb_inst_5_douta[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_183 (
  .O(mux_o_183),
  .I0(dpb_inst_6_douta[12]),
  .I1(dpb_inst_7_douta[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(dpb_inst_8_douta[12]),
  .I1(dpb_inst_9_douta[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_185 (
  .O(mux_o_185),
  .I0(dpb_inst_10_douta[12]),
  .I1(dpb_inst_11_douta[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_186 (
  .O(mux_o_186),
  .I0(dpb_inst_12_douta[12]),
  .I1(dpb_inst_13_douta[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_187 (
  .O(mux_o_187),
  .I0(dpb_inst_14_douta[12]),
  .I1(dpb_inst_15_douta[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_188 (
  .O(mux_o_188),
  .I0(mux_o_180),
  .I1(mux_o_181),
  .S0(dff_q_2)
);
MUX2 mux_inst_189 (
  .O(mux_o_189),
  .I0(mux_o_182),
  .I1(mux_o_183),
  .S0(dff_q_2)
);
MUX2 mux_inst_190 (
  .O(mux_o_190),
  .I0(mux_o_184),
  .I1(mux_o_185),
  .S0(dff_q_2)
);
MUX2 mux_inst_191 (
  .O(mux_o_191),
  .I0(mux_o_186),
  .I1(mux_o_187),
  .S0(dff_q_2)
);
MUX2 mux_inst_192 (
  .O(mux_o_192),
  .I0(mux_o_188),
  .I1(mux_o_189),
  .S0(dff_q_1)
);
MUX2 mux_inst_193 (
  .O(mux_o_193),
  .I0(mux_o_190),
  .I1(mux_o_191),
  .S0(dff_q_1)
);
MUX2 mux_inst_194 (
  .O(douta[12]),
  .I0(mux_o_192),
  .I1(mux_o_193),
  .S0(dff_q_0)
);
MUX2 mux_inst_195 (
  .O(mux_o_195),
  .I0(dpb_inst_0_douta[13]),
  .I1(dpb_inst_1_douta[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_196 (
  .O(mux_o_196),
  .I0(dpb_inst_2_douta[13]),
  .I1(dpb_inst_3_douta[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_197 (
  .O(mux_o_197),
  .I0(dpb_inst_4_douta[13]),
  .I1(dpb_inst_5_douta[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_198 (
  .O(mux_o_198),
  .I0(dpb_inst_6_douta[13]),
  .I1(dpb_inst_7_douta[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_199 (
  .O(mux_o_199),
  .I0(dpb_inst_8_douta[13]),
  .I1(dpb_inst_9_douta[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_200 (
  .O(mux_o_200),
  .I0(dpb_inst_10_douta[13]),
  .I1(dpb_inst_11_douta[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_201 (
  .O(mux_o_201),
  .I0(dpb_inst_12_douta[13]),
  .I1(dpb_inst_13_douta[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_202 (
  .O(mux_o_202),
  .I0(dpb_inst_14_douta[13]),
  .I1(dpb_inst_15_douta[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_203 (
  .O(mux_o_203),
  .I0(mux_o_195),
  .I1(mux_o_196),
  .S0(dff_q_2)
);
MUX2 mux_inst_204 (
  .O(mux_o_204),
  .I0(mux_o_197),
  .I1(mux_o_198),
  .S0(dff_q_2)
);
MUX2 mux_inst_205 (
  .O(mux_o_205),
  .I0(mux_o_199),
  .I1(mux_o_200),
  .S0(dff_q_2)
);
MUX2 mux_inst_206 (
  .O(mux_o_206),
  .I0(mux_o_201),
  .I1(mux_o_202),
  .S0(dff_q_2)
);
MUX2 mux_inst_207 (
  .O(mux_o_207),
  .I0(mux_o_203),
  .I1(mux_o_204),
  .S0(dff_q_1)
);
MUX2 mux_inst_208 (
  .O(mux_o_208),
  .I0(mux_o_205),
  .I1(mux_o_206),
  .S0(dff_q_1)
);
MUX2 mux_inst_209 (
  .O(douta[13]),
  .I0(mux_o_207),
  .I1(mux_o_208),
  .S0(dff_q_0)
);
MUX2 mux_inst_210 (
  .O(mux_o_210),
  .I0(dpb_inst_0_douta[14]),
  .I1(dpb_inst_1_douta[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_211 (
  .O(mux_o_211),
  .I0(dpb_inst_2_douta[14]),
  .I1(dpb_inst_3_douta[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_212 (
  .O(mux_o_212),
  .I0(dpb_inst_4_douta[14]),
  .I1(dpb_inst_5_douta[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_213 (
  .O(mux_o_213),
  .I0(dpb_inst_6_douta[14]),
  .I1(dpb_inst_7_douta[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_214 (
  .O(mux_o_214),
  .I0(dpb_inst_8_douta[14]),
  .I1(dpb_inst_9_douta[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_215 (
  .O(mux_o_215),
  .I0(dpb_inst_10_douta[14]),
  .I1(dpb_inst_11_douta[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_216 (
  .O(mux_o_216),
  .I0(dpb_inst_12_douta[14]),
  .I1(dpb_inst_13_douta[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_217 (
  .O(mux_o_217),
  .I0(dpb_inst_14_douta[14]),
  .I1(dpb_inst_15_douta[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_218 (
  .O(mux_o_218),
  .I0(mux_o_210),
  .I1(mux_o_211),
  .S0(dff_q_2)
);
MUX2 mux_inst_219 (
  .O(mux_o_219),
  .I0(mux_o_212),
  .I1(mux_o_213),
  .S0(dff_q_2)
);
MUX2 mux_inst_220 (
  .O(mux_o_220),
  .I0(mux_o_214),
  .I1(mux_o_215),
  .S0(dff_q_2)
);
MUX2 mux_inst_221 (
  .O(mux_o_221),
  .I0(mux_o_216),
  .I1(mux_o_217),
  .S0(dff_q_2)
);
MUX2 mux_inst_222 (
  .O(mux_o_222),
  .I0(mux_o_218),
  .I1(mux_o_219),
  .S0(dff_q_1)
);
MUX2 mux_inst_223 (
  .O(mux_o_223),
  .I0(mux_o_220),
  .I1(mux_o_221),
  .S0(dff_q_1)
);
MUX2 mux_inst_224 (
  .O(douta[14]),
  .I0(mux_o_222),
  .I1(mux_o_223),
  .S0(dff_q_0)
);
MUX2 mux_inst_225 (
  .O(mux_o_225),
  .I0(dpb_inst_0_douta[15]),
  .I1(dpb_inst_1_douta[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_226 (
  .O(mux_o_226),
  .I0(dpb_inst_2_douta[15]),
  .I1(dpb_inst_3_douta[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_227 (
  .O(mux_o_227),
  .I0(dpb_inst_4_douta[15]),
  .I1(dpb_inst_5_douta[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_228 (
  .O(mux_o_228),
  .I0(dpb_inst_6_douta[15]),
  .I1(dpb_inst_7_douta[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_229 (
  .O(mux_o_229),
  .I0(dpb_inst_8_douta[15]),
  .I1(dpb_inst_9_douta[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_230 (
  .O(mux_o_230),
  .I0(dpb_inst_10_douta[15]),
  .I1(dpb_inst_11_douta[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_231 (
  .O(mux_o_231),
  .I0(dpb_inst_12_douta[15]),
  .I1(dpb_inst_13_douta[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_232 (
  .O(mux_o_232),
  .I0(dpb_inst_14_douta[15]),
  .I1(dpb_inst_15_douta[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_233 (
  .O(mux_o_233),
  .I0(mux_o_225),
  .I1(mux_o_226),
  .S0(dff_q_2)
);
MUX2 mux_inst_234 (
  .O(mux_o_234),
  .I0(mux_o_227),
  .I1(mux_o_228),
  .S0(dff_q_2)
);
MUX2 mux_inst_235 (
  .O(mux_o_235),
  .I0(mux_o_229),
  .I1(mux_o_230),
  .S0(dff_q_2)
);
MUX2 mux_inst_236 (
  .O(mux_o_236),
  .I0(mux_o_231),
  .I1(mux_o_232),
  .S0(dff_q_2)
);
MUX2 mux_inst_237 (
  .O(mux_o_237),
  .I0(mux_o_233),
  .I1(mux_o_234),
  .S0(dff_q_1)
);
MUX2 mux_inst_238 (
  .O(mux_o_238),
  .I0(mux_o_235),
  .I1(mux_o_236),
  .S0(dff_q_1)
);
MUX2 mux_inst_239 (
  .O(douta[15]),
  .I0(mux_o_237),
  .I1(mux_o_238),
  .S0(dff_q_0)
);
MUX2 mux_inst_240 (
  .O(mux_o_240),
  .I0(dpb_inst_16_douta[16]),
  .I1(dpb_inst_17_douta[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_241 (
  .O(mux_o_241),
  .I0(dpb_inst_18_douta[16]),
  .I1(dpb_inst_19_douta[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_242 (
  .O(mux_o_242),
  .I0(dpb_inst_20_douta[16]),
  .I1(dpb_inst_21_douta[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_243 (
  .O(mux_o_243),
  .I0(dpb_inst_22_douta[16]),
  .I1(dpb_inst_23_douta[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_244 (
  .O(mux_o_244),
  .I0(dpb_inst_24_douta[16]),
  .I1(dpb_inst_25_douta[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_245 (
  .O(mux_o_245),
  .I0(dpb_inst_26_douta[16]),
  .I1(dpb_inst_27_douta[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_246 (
  .O(mux_o_246),
  .I0(dpb_inst_28_douta[16]),
  .I1(dpb_inst_29_douta[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_247 (
  .O(mux_o_247),
  .I0(dpb_inst_30_douta[16]),
  .I1(dpb_inst_31_douta[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_248 (
  .O(mux_o_248),
  .I0(mux_o_240),
  .I1(mux_o_241),
  .S0(dff_q_2)
);
MUX2 mux_inst_249 (
  .O(mux_o_249),
  .I0(mux_o_242),
  .I1(mux_o_243),
  .S0(dff_q_2)
);
MUX2 mux_inst_250 (
  .O(mux_o_250),
  .I0(mux_o_244),
  .I1(mux_o_245),
  .S0(dff_q_2)
);
MUX2 mux_inst_251 (
  .O(mux_o_251),
  .I0(mux_o_246),
  .I1(mux_o_247),
  .S0(dff_q_2)
);
MUX2 mux_inst_252 (
  .O(mux_o_252),
  .I0(mux_o_248),
  .I1(mux_o_249),
  .S0(dff_q_1)
);
MUX2 mux_inst_253 (
  .O(mux_o_253),
  .I0(mux_o_250),
  .I1(mux_o_251),
  .S0(dff_q_1)
);
MUX2 mux_inst_254 (
  .O(douta[16]),
  .I0(mux_o_252),
  .I1(mux_o_253),
  .S0(dff_q_0)
);
MUX2 mux_inst_255 (
  .O(mux_o_255),
  .I0(dpb_inst_16_douta[17]),
  .I1(dpb_inst_17_douta[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_256 (
  .O(mux_o_256),
  .I0(dpb_inst_18_douta[17]),
  .I1(dpb_inst_19_douta[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_257 (
  .O(mux_o_257),
  .I0(dpb_inst_20_douta[17]),
  .I1(dpb_inst_21_douta[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_258 (
  .O(mux_o_258),
  .I0(dpb_inst_22_douta[17]),
  .I1(dpb_inst_23_douta[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_259 (
  .O(mux_o_259),
  .I0(dpb_inst_24_douta[17]),
  .I1(dpb_inst_25_douta[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_260 (
  .O(mux_o_260),
  .I0(dpb_inst_26_douta[17]),
  .I1(dpb_inst_27_douta[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_261 (
  .O(mux_o_261),
  .I0(dpb_inst_28_douta[17]),
  .I1(dpb_inst_29_douta[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_262 (
  .O(mux_o_262),
  .I0(dpb_inst_30_douta[17]),
  .I1(dpb_inst_31_douta[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_263 (
  .O(mux_o_263),
  .I0(mux_o_255),
  .I1(mux_o_256),
  .S0(dff_q_2)
);
MUX2 mux_inst_264 (
  .O(mux_o_264),
  .I0(mux_o_257),
  .I1(mux_o_258),
  .S0(dff_q_2)
);
MUX2 mux_inst_265 (
  .O(mux_o_265),
  .I0(mux_o_259),
  .I1(mux_o_260),
  .S0(dff_q_2)
);
MUX2 mux_inst_266 (
  .O(mux_o_266),
  .I0(mux_o_261),
  .I1(mux_o_262),
  .S0(dff_q_2)
);
MUX2 mux_inst_267 (
  .O(mux_o_267),
  .I0(mux_o_263),
  .I1(mux_o_264),
  .S0(dff_q_1)
);
MUX2 mux_inst_268 (
  .O(mux_o_268),
  .I0(mux_o_265),
  .I1(mux_o_266),
  .S0(dff_q_1)
);
MUX2 mux_inst_269 (
  .O(douta[17]),
  .I0(mux_o_267),
  .I1(mux_o_268),
  .S0(dff_q_0)
);
MUX2 mux_inst_270 (
  .O(mux_o_270),
  .I0(dpb_inst_16_douta[18]),
  .I1(dpb_inst_17_douta[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_271 (
  .O(mux_o_271),
  .I0(dpb_inst_18_douta[18]),
  .I1(dpb_inst_19_douta[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_272 (
  .O(mux_o_272),
  .I0(dpb_inst_20_douta[18]),
  .I1(dpb_inst_21_douta[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_273 (
  .O(mux_o_273),
  .I0(dpb_inst_22_douta[18]),
  .I1(dpb_inst_23_douta[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_274 (
  .O(mux_o_274),
  .I0(dpb_inst_24_douta[18]),
  .I1(dpb_inst_25_douta[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_275 (
  .O(mux_o_275),
  .I0(dpb_inst_26_douta[18]),
  .I1(dpb_inst_27_douta[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_276 (
  .O(mux_o_276),
  .I0(dpb_inst_28_douta[18]),
  .I1(dpb_inst_29_douta[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_277 (
  .O(mux_o_277),
  .I0(dpb_inst_30_douta[18]),
  .I1(dpb_inst_31_douta[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_278 (
  .O(mux_o_278),
  .I0(mux_o_270),
  .I1(mux_o_271),
  .S0(dff_q_2)
);
MUX2 mux_inst_279 (
  .O(mux_o_279),
  .I0(mux_o_272),
  .I1(mux_o_273),
  .S0(dff_q_2)
);
MUX2 mux_inst_280 (
  .O(mux_o_280),
  .I0(mux_o_274),
  .I1(mux_o_275),
  .S0(dff_q_2)
);
MUX2 mux_inst_281 (
  .O(mux_o_281),
  .I0(mux_o_276),
  .I1(mux_o_277),
  .S0(dff_q_2)
);
MUX2 mux_inst_282 (
  .O(mux_o_282),
  .I0(mux_o_278),
  .I1(mux_o_279),
  .S0(dff_q_1)
);
MUX2 mux_inst_283 (
  .O(mux_o_283),
  .I0(mux_o_280),
  .I1(mux_o_281),
  .S0(dff_q_1)
);
MUX2 mux_inst_284 (
  .O(douta[18]),
  .I0(mux_o_282),
  .I1(mux_o_283),
  .S0(dff_q_0)
);
MUX2 mux_inst_285 (
  .O(mux_o_285),
  .I0(dpb_inst_16_douta[19]),
  .I1(dpb_inst_17_douta[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_286 (
  .O(mux_o_286),
  .I0(dpb_inst_18_douta[19]),
  .I1(dpb_inst_19_douta[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_287 (
  .O(mux_o_287),
  .I0(dpb_inst_20_douta[19]),
  .I1(dpb_inst_21_douta[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_288 (
  .O(mux_o_288),
  .I0(dpb_inst_22_douta[19]),
  .I1(dpb_inst_23_douta[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_289 (
  .O(mux_o_289),
  .I0(dpb_inst_24_douta[19]),
  .I1(dpb_inst_25_douta[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_290 (
  .O(mux_o_290),
  .I0(dpb_inst_26_douta[19]),
  .I1(dpb_inst_27_douta[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_291 (
  .O(mux_o_291),
  .I0(dpb_inst_28_douta[19]),
  .I1(dpb_inst_29_douta[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_292 (
  .O(mux_o_292),
  .I0(dpb_inst_30_douta[19]),
  .I1(dpb_inst_31_douta[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_293 (
  .O(mux_o_293),
  .I0(mux_o_285),
  .I1(mux_o_286),
  .S0(dff_q_2)
);
MUX2 mux_inst_294 (
  .O(mux_o_294),
  .I0(mux_o_287),
  .I1(mux_o_288),
  .S0(dff_q_2)
);
MUX2 mux_inst_295 (
  .O(mux_o_295),
  .I0(mux_o_289),
  .I1(mux_o_290),
  .S0(dff_q_2)
);
MUX2 mux_inst_296 (
  .O(mux_o_296),
  .I0(mux_o_291),
  .I1(mux_o_292),
  .S0(dff_q_2)
);
MUX2 mux_inst_297 (
  .O(mux_o_297),
  .I0(mux_o_293),
  .I1(mux_o_294),
  .S0(dff_q_1)
);
MUX2 mux_inst_298 (
  .O(mux_o_298),
  .I0(mux_o_295),
  .I1(mux_o_296),
  .S0(dff_q_1)
);
MUX2 mux_inst_299 (
  .O(douta[19]),
  .I0(mux_o_297),
  .I1(mux_o_298),
  .S0(dff_q_0)
);
MUX2 mux_inst_300 (
  .O(mux_o_300),
  .I0(dpb_inst_16_douta[20]),
  .I1(dpb_inst_17_douta[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_301 (
  .O(mux_o_301),
  .I0(dpb_inst_18_douta[20]),
  .I1(dpb_inst_19_douta[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_302 (
  .O(mux_o_302),
  .I0(dpb_inst_20_douta[20]),
  .I1(dpb_inst_21_douta[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_303 (
  .O(mux_o_303),
  .I0(dpb_inst_22_douta[20]),
  .I1(dpb_inst_23_douta[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_304 (
  .O(mux_o_304),
  .I0(dpb_inst_24_douta[20]),
  .I1(dpb_inst_25_douta[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_305 (
  .O(mux_o_305),
  .I0(dpb_inst_26_douta[20]),
  .I1(dpb_inst_27_douta[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_306 (
  .O(mux_o_306),
  .I0(dpb_inst_28_douta[20]),
  .I1(dpb_inst_29_douta[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_307 (
  .O(mux_o_307),
  .I0(dpb_inst_30_douta[20]),
  .I1(dpb_inst_31_douta[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_308 (
  .O(mux_o_308),
  .I0(mux_o_300),
  .I1(mux_o_301),
  .S0(dff_q_2)
);
MUX2 mux_inst_309 (
  .O(mux_o_309),
  .I0(mux_o_302),
  .I1(mux_o_303),
  .S0(dff_q_2)
);
MUX2 mux_inst_310 (
  .O(mux_o_310),
  .I0(mux_o_304),
  .I1(mux_o_305),
  .S0(dff_q_2)
);
MUX2 mux_inst_311 (
  .O(mux_o_311),
  .I0(mux_o_306),
  .I1(mux_o_307),
  .S0(dff_q_2)
);
MUX2 mux_inst_312 (
  .O(mux_o_312),
  .I0(mux_o_308),
  .I1(mux_o_309),
  .S0(dff_q_1)
);
MUX2 mux_inst_313 (
  .O(mux_o_313),
  .I0(mux_o_310),
  .I1(mux_o_311),
  .S0(dff_q_1)
);
MUX2 mux_inst_314 (
  .O(douta[20]),
  .I0(mux_o_312),
  .I1(mux_o_313),
  .S0(dff_q_0)
);
MUX2 mux_inst_315 (
  .O(mux_o_315),
  .I0(dpb_inst_16_douta[21]),
  .I1(dpb_inst_17_douta[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_316 (
  .O(mux_o_316),
  .I0(dpb_inst_18_douta[21]),
  .I1(dpb_inst_19_douta[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_317 (
  .O(mux_o_317),
  .I0(dpb_inst_20_douta[21]),
  .I1(dpb_inst_21_douta[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_318 (
  .O(mux_o_318),
  .I0(dpb_inst_22_douta[21]),
  .I1(dpb_inst_23_douta[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_319 (
  .O(mux_o_319),
  .I0(dpb_inst_24_douta[21]),
  .I1(dpb_inst_25_douta[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_320 (
  .O(mux_o_320),
  .I0(dpb_inst_26_douta[21]),
  .I1(dpb_inst_27_douta[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_321 (
  .O(mux_o_321),
  .I0(dpb_inst_28_douta[21]),
  .I1(dpb_inst_29_douta[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_322 (
  .O(mux_o_322),
  .I0(dpb_inst_30_douta[21]),
  .I1(dpb_inst_31_douta[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_323 (
  .O(mux_o_323),
  .I0(mux_o_315),
  .I1(mux_o_316),
  .S0(dff_q_2)
);
MUX2 mux_inst_324 (
  .O(mux_o_324),
  .I0(mux_o_317),
  .I1(mux_o_318),
  .S0(dff_q_2)
);
MUX2 mux_inst_325 (
  .O(mux_o_325),
  .I0(mux_o_319),
  .I1(mux_o_320),
  .S0(dff_q_2)
);
MUX2 mux_inst_326 (
  .O(mux_o_326),
  .I0(mux_o_321),
  .I1(mux_o_322),
  .S0(dff_q_2)
);
MUX2 mux_inst_327 (
  .O(mux_o_327),
  .I0(mux_o_323),
  .I1(mux_o_324),
  .S0(dff_q_1)
);
MUX2 mux_inst_328 (
  .O(mux_o_328),
  .I0(mux_o_325),
  .I1(mux_o_326),
  .S0(dff_q_1)
);
MUX2 mux_inst_329 (
  .O(douta[21]),
  .I0(mux_o_327),
  .I1(mux_o_328),
  .S0(dff_q_0)
);
MUX2 mux_inst_330 (
  .O(mux_o_330),
  .I0(dpb_inst_16_douta[22]),
  .I1(dpb_inst_17_douta[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_331 (
  .O(mux_o_331),
  .I0(dpb_inst_18_douta[22]),
  .I1(dpb_inst_19_douta[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_332 (
  .O(mux_o_332),
  .I0(dpb_inst_20_douta[22]),
  .I1(dpb_inst_21_douta[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_333 (
  .O(mux_o_333),
  .I0(dpb_inst_22_douta[22]),
  .I1(dpb_inst_23_douta[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_334 (
  .O(mux_o_334),
  .I0(dpb_inst_24_douta[22]),
  .I1(dpb_inst_25_douta[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_335 (
  .O(mux_o_335),
  .I0(dpb_inst_26_douta[22]),
  .I1(dpb_inst_27_douta[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_336 (
  .O(mux_o_336),
  .I0(dpb_inst_28_douta[22]),
  .I1(dpb_inst_29_douta[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_337 (
  .O(mux_o_337),
  .I0(dpb_inst_30_douta[22]),
  .I1(dpb_inst_31_douta[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_338 (
  .O(mux_o_338),
  .I0(mux_o_330),
  .I1(mux_o_331),
  .S0(dff_q_2)
);
MUX2 mux_inst_339 (
  .O(mux_o_339),
  .I0(mux_o_332),
  .I1(mux_o_333),
  .S0(dff_q_2)
);
MUX2 mux_inst_340 (
  .O(mux_o_340),
  .I0(mux_o_334),
  .I1(mux_o_335),
  .S0(dff_q_2)
);
MUX2 mux_inst_341 (
  .O(mux_o_341),
  .I0(mux_o_336),
  .I1(mux_o_337),
  .S0(dff_q_2)
);
MUX2 mux_inst_342 (
  .O(mux_o_342),
  .I0(mux_o_338),
  .I1(mux_o_339),
  .S0(dff_q_1)
);
MUX2 mux_inst_343 (
  .O(mux_o_343),
  .I0(mux_o_340),
  .I1(mux_o_341),
  .S0(dff_q_1)
);
MUX2 mux_inst_344 (
  .O(douta[22]),
  .I0(mux_o_342),
  .I1(mux_o_343),
  .S0(dff_q_0)
);
MUX2 mux_inst_345 (
  .O(mux_o_345),
  .I0(dpb_inst_16_douta[23]),
  .I1(dpb_inst_17_douta[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_346 (
  .O(mux_o_346),
  .I0(dpb_inst_18_douta[23]),
  .I1(dpb_inst_19_douta[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_347 (
  .O(mux_o_347),
  .I0(dpb_inst_20_douta[23]),
  .I1(dpb_inst_21_douta[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_348 (
  .O(mux_o_348),
  .I0(dpb_inst_22_douta[23]),
  .I1(dpb_inst_23_douta[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_349 (
  .O(mux_o_349),
  .I0(dpb_inst_24_douta[23]),
  .I1(dpb_inst_25_douta[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_350 (
  .O(mux_o_350),
  .I0(dpb_inst_26_douta[23]),
  .I1(dpb_inst_27_douta[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_351 (
  .O(mux_o_351),
  .I0(dpb_inst_28_douta[23]),
  .I1(dpb_inst_29_douta[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_352 (
  .O(mux_o_352),
  .I0(dpb_inst_30_douta[23]),
  .I1(dpb_inst_31_douta[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_353 (
  .O(mux_o_353),
  .I0(mux_o_345),
  .I1(mux_o_346),
  .S0(dff_q_2)
);
MUX2 mux_inst_354 (
  .O(mux_o_354),
  .I0(mux_o_347),
  .I1(mux_o_348),
  .S0(dff_q_2)
);
MUX2 mux_inst_355 (
  .O(mux_o_355),
  .I0(mux_o_349),
  .I1(mux_o_350),
  .S0(dff_q_2)
);
MUX2 mux_inst_356 (
  .O(mux_o_356),
  .I0(mux_o_351),
  .I1(mux_o_352),
  .S0(dff_q_2)
);
MUX2 mux_inst_357 (
  .O(mux_o_357),
  .I0(mux_o_353),
  .I1(mux_o_354),
  .S0(dff_q_1)
);
MUX2 mux_inst_358 (
  .O(mux_o_358),
  .I0(mux_o_355),
  .I1(mux_o_356),
  .S0(dff_q_1)
);
MUX2 mux_inst_359 (
  .O(douta[23]),
  .I0(mux_o_357),
  .I1(mux_o_358),
  .S0(dff_q_0)
);
MUX2 mux_inst_360 (
  .O(mux_o_360),
  .I0(dpb_inst_16_douta[24]),
  .I1(dpb_inst_17_douta[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_361 (
  .O(mux_o_361),
  .I0(dpb_inst_18_douta[24]),
  .I1(dpb_inst_19_douta[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_362 (
  .O(mux_o_362),
  .I0(dpb_inst_20_douta[24]),
  .I1(dpb_inst_21_douta[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_363 (
  .O(mux_o_363),
  .I0(dpb_inst_22_douta[24]),
  .I1(dpb_inst_23_douta[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_364 (
  .O(mux_o_364),
  .I0(dpb_inst_24_douta[24]),
  .I1(dpb_inst_25_douta[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_365 (
  .O(mux_o_365),
  .I0(dpb_inst_26_douta[24]),
  .I1(dpb_inst_27_douta[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_366 (
  .O(mux_o_366),
  .I0(dpb_inst_28_douta[24]),
  .I1(dpb_inst_29_douta[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_367 (
  .O(mux_o_367),
  .I0(dpb_inst_30_douta[24]),
  .I1(dpb_inst_31_douta[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_368 (
  .O(mux_o_368),
  .I0(mux_o_360),
  .I1(mux_o_361),
  .S0(dff_q_2)
);
MUX2 mux_inst_369 (
  .O(mux_o_369),
  .I0(mux_o_362),
  .I1(mux_o_363),
  .S0(dff_q_2)
);
MUX2 mux_inst_370 (
  .O(mux_o_370),
  .I0(mux_o_364),
  .I1(mux_o_365),
  .S0(dff_q_2)
);
MUX2 mux_inst_371 (
  .O(mux_o_371),
  .I0(mux_o_366),
  .I1(mux_o_367),
  .S0(dff_q_2)
);
MUX2 mux_inst_372 (
  .O(mux_o_372),
  .I0(mux_o_368),
  .I1(mux_o_369),
  .S0(dff_q_1)
);
MUX2 mux_inst_373 (
  .O(mux_o_373),
  .I0(mux_o_370),
  .I1(mux_o_371),
  .S0(dff_q_1)
);
MUX2 mux_inst_374 (
  .O(douta[24]),
  .I0(mux_o_372),
  .I1(mux_o_373),
  .S0(dff_q_0)
);
MUX2 mux_inst_375 (
  .O(mux_o_375),
  .I0(dpb_inst_16_douta[25]),
  .I1(dpb_inst_17_douta[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_376 (
  .O(mux_o_376),
  .I0(dpb_inst_18_douta[25]),
  .I1(dpb_inst_19_douta[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_377 (
  .O(mux_o_377),
  .I0(dpb_inst_20_douta[25]),
  .I1(dpb_inst_21_douta[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_378 (
  .O(mux_o_378),
  .I0(dpb_inst_22_douta[25]),
  .I1(dpb_inst_23_douta[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_379 (
  .O(mux_o_379),
  .I0(dpb_inst_24_douta[25]),
  .I1(dpb_inst_25_douta[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_380 (
  .O(mux_o_380),
  .I0(dpb_inst_26_douta[25]),
  .I1(dpb_inst_27_douta[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_381 (
  .O(mux_o_381),
  .I0(dpb_inst_28_douta[25]),
  .I1(dpb_inst_29_douta[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_382 (
  .O(mux_o_382),
  .I0(dpb_inst_30_douta[25]),
  .I1(dpb_inst_31_douta[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_383 (
  .O(mux_o_383),
  .I0(mux_o_375),
  .I1(mux_o_376),
  .S0(dff_q_2)
);
MUX2 mux_inst_384 (
  .O(mux_o_384),
  .I0(mux_o_377),
  .I1(mux_o_378),
  .S0(dff_q_2)
);
MUX2 mux_inst_385 (
  .O(mux_o_385),
  .I0(mux_o_379),
  .I1(mux_o_380),
  .S0(dff_q_2)
);
MUX2 mux_inst_386 (
  .O(mux_o_386),
  .I0(mux_o_381),
  .I1(mux_o_382),
  .S0(dff_q_2)
);
MUX2 mux_inst_387 (
  .O(mux_o_387),
  .I0(mux_o_383),
  .I1(mux_o_384),
  .S0(dff_q_1)
);
MUX2 mux_inst_388 (
  .O(mux_o_388),
  .I0(mux_o_385),
  .I1(mux_o_386),
  .S0(dff_q_1)
);
MUX2 mux_inst_389 (
  .O(douta[25]),
  .I0(mux_o_387),
  .I1(mux_o_388),
  .S0(dff_q_0)
);
MUX2 mux_inst_390 (
  .O(mux_o_390),
  .I0(dpb_inst_16_douta[26]),
  .I1(dpb_inst_17_douta[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_391 (
  .O(mux_o_391),
  .I0(dpb_inst_18_douta[26]),
  .I1(dpb_inst_19_douta[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_392 (
  .O(mux_o_392),
  .I0(dpb_inst_20_douta[26]),
  .I1(dpb_inst_21_douta[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_393 (
  .O(mux_o_393),
  .I0(dpb_inst_22_douta[26]),
  .I1(dpb_inst_23_douta[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_394 (
  .O(mux_o_394),
  .I0(dpb_inst_24_douta[26]),
  .I1(dpb_inst_25_douta[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_395 (
  .O(mux_o_395),
  .I0(dpb_inst_26_douta[26]),
  .I1(dpb_inst_27_douta[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_396 (
  .O(mux_o_396),
  .I0(dpb_inst_28_douta[26]),
  .I1(dpb_inst_29_douta[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_397 (
  .O(mux_o_397),
  .I0(dpb_inst_30_douta[26]),
  .I1(dpb_inst_31_douta[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_398 (
  .O(mux_o_398),
  .I0(mux_o_390),
  .I1(mux_o_391),
  .S0(dff_q_2)
);
MUX2 mux_inst_399 (
  .O(mux_o_399),
  .I0(mux_o_392),
  .I1(mux_o_393),
  .S0(dff_q_2)
);
MUX2 mux_inst_400 (
  .O(mux_o_400),
  .I0(mux_o_394),
  .I1(mux_o_395),
  .S0(dff_q_2)
);
MUX2 mux_inst_401 (
  .O(mux_o_401),
  .I0(mux_o_396),
  .I1(mux_o_397),
  .S0(dff_q_2)
);
MUX2 mux_inst_402 (
  .O(mux_o_402),
  .I0(mux_o_398),
  .I1(mux_o_399),
  .S0(dff_q_1)
);
MUX2 mux_inst_403 (
  .O(mux_o_403),
  .I0(mux_o_400),
  .I1(mux_o_401),
  .S0(dff_q_1)
);
MUX2 mux_inst_404 (
  .O(douta[26]),
  .I0(mux_o_402),
  .I1(mux_o_403),
  .S0(dff_q_0)
);
MUX2 mux_inst_405 (
  .O(mux_o_405),
  .I0(dpb_inst_16_douta[27]),
  .I1(dpb_inst_17_douta[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_406 (
  .O(mux_o_406),
  .I0(dpb_inst_18_douta[27]),
  .I1(dpb_inst_19_douta[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_407 (
  .O(mux_o_407),
  .I0(dpb_inst_20_douta[27]),
  .I1(dpb_inst_21_douta[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_408 (
  .O(mux_o_408),
  .I0(dpb_inst_22_douta[27]),
  .I1(dpb_inst_23_douta[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_409 (
  .O(mux_o_409),
  .I0(dpb_inst_24_douta[27]),
  .I1(dpb_inst_25_douta[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_410 (
  .O(mux_o_410),
  .I0(dpb_inst_26_douta[27]),
  .I1(dpb_inst_27_douta[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_411 (
  .O(mux_o_411),
  .I0(dpb_inst_28_douta[27]),
  .I1(dpb_inst_29_douta[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_412 (
  .O(mux_o_412),
  .I0(dpb_inst_30_douta[27]),
  .I1(dpb_inst_31_douta[27]),
  .S0(dff_q_3)
);
MUX2 mux_inst_413 (
  .O(mux_o_413),
  .I0(mux_o_405),
  .I1(mux_o_406),
  .S0(dff_q_2)
);
MUX2 mux_inst_414 (
  .O(mux_o_414),
  .I0(mux_o_407),
  .I1(mux_o_408),
  .S0(dff_q_2)
);
MUX2 mux_inst_415 (
  .O(mux_o_415),
  .I0(mux_o_409),
  .I1(mux_o_410),
  .S0(dff_q_2)
);
MUX2 mux_inst_416 (
  .O(mux_o_416),
  .I0(mux_o_411),
  .I1(mux_o_412),
  .S0(dff_q_2)
);
MUX2 mux_inst_417 (
  .O(mux_o_417),
  .I0(mux_o_413),
  .I1(mux_o_414),
  .S0(dff_q_1)
);
MUX2 mux_inst_418 (
  .O(mux_o_418),
  .I0(mux_o_415),
  .I1(mux_o_416),
  .S0(dff_q_1)
);
MUX2 mux_inst_419 (
  .O(douta[27]),
  .I0(mux_o_417),
  .I1(mux_o_418),
  .S0(dff_q_0)
);
MUX2 mux_inst_420 (
  .O(mux_o_420),
  .I0(dpb_inst_16_douta[28]),
  .I1(dpb_inst_17_douta[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_421 (
  .O(mux_o_421),
  .I0(dpb_inst_18_douta[28]),
  .I1(dpb_inst_19_douta[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_422 (
  .O(mux_o_422),
  .I0(dpb_inst_20_douta[28]),
  .I1(dpb_inst_21_douta[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_423 (
  .O(mux_o_423),
  .I0(dpb_inst_22_douta[28]),
  .I1(dpb_inst_23_douta[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_424 (
  .O(mux_o_424),
  .I0(dpb_inst_24_douta[28]),
  .I1(dpb_inst_25_douta[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_425 (
  .O(mux_o_425),
  .I0(dpb_inst_26_douta[28]),
  .I1(dpb_inst_27_douta[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_426 (
  .O(mux_o_426),
  .I0(dpb_inst_28_douta[28]),
  .I1(dpb_inst_29_douta[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_427 (
  .O(mux_o_427),
  .I0(dpb_inst_30_douta[28]),
  .I1(dpb_inst_31_douta[28]),
  .S0(dff_q_3)
);
MUX2 mux_inst_428 (
  .O(mux_o_428),
  .I0(mux_o_420),
  .I1(mux_o_421),
  .S0(dff_q_2)
);
MUX2 mux_inst_429 (
  .O(mux_o_429),
  .I0(mux_o_422),
  .I1(mux_o_423),
  .S0(dff_q_2)
);
MUX2 mux_inst_430 (
  .O(mux_o_430),
  .I0(mux_o_424),
  .I1(mux_o_425),
  .S0(dff_q_2)
);
MUX2 mux_inst_431 (
  .O(mux_o_431),
  .I0(mux_o_426),
  .I1(mux_o_427),
  .S0(dff_q_2)
);
MUX2 mux_inst_432 (
  .O(mux_o_432),
  .I0(mux_o_428),
  .I1(mux_o_429),
  .S0(dff_q_1)
);
MUX2 mux_inst_433 (
  .O(mux_o_433),
  .I0(mux_o_430),
  .I1(mux_o_431),
  .S0(dff_q_1)
);
MUX2 mux_inst_434 (
  .O(douta[28]),
  .I0(mux_o_432),
  .I1(mux_o_433),
  .S0(dff_q_0)
);
MUX2 mux_inst_435 (
  .O(mux_o_435),
  .I0(dpb_inst_16_douta[29]),
  .I1(dpb_inst_17_douta[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_436 (
  .O(mux_o_436),
  .I0(dpb_inst_18_douta[29]),
  .I1(dpb_inst_19_douta[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_437 (
  .O(mux_o_437),
  .I0(dpb_inst_20_douta[29]),
  .I1(dpb_inst_21_douta[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_438 (
  .O(mux_o_438),
  .I0(dpb_inst_22_douta[29]),
  .I1(dpb_inst_23_douta[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_439 (
  .O(mux_o_439),
  .I0(dpb_inst_24_douta[29]),
  .I1(dpb_inst_25_douta[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_440 (
  .O(mux_o_440),
  .I0(dpb_inst_26_douta[29]),
  .I1(dpb_inst_27_douta[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_441 (
  .O(mux_o_441),
  .I0(dpb_inst_28_douta[29]),
  .I1(dpb_inst_29_douta[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_442 (
  .O(mux_o_442),
  .I0(dpb_inst_30_douta[29]),
  .I1(dpb_inst_31_douta[29]),
  .S0(dff_q_3)
);
MUX2 mux_inst_443 (
  .O(mux_o_443),
  .I0(mux_o_435),
  .I1(mux_o_436),
  .S0(dff_q_2)
);
MUX2 mux_inst_444 (
  .O(mux_o_444),
  .I0(mux_o_437),
  .I1(mux_o_438),
  .S0(dff_q_2)
);
MUX2 mux_inst_445 (
  .O(mux_o_445),
  .I0(mux_o_439),
  .I1(mux_o_440),
  .S0(dff_q_2)
);
MUX2 mux_inst_446 (
  .O(mux_o_446),
  .I0(mux_o_441),
  .I1(mux_o_442),
  .S0(dff_q_2)
);
MUX2 mux_inst_447 (
  .O(mux_o_447),
  .I0(mux_o_443),
  .I1(mux_o_444),
  .S0(dff_q_1)
);
MUX2 mux_inst_448 (
  .O(mux_o_448),
  .I0(mux_o_445),
  .I1(mux_o_446),
  .S0(dff_q_1)
);
MUX2 mux_inst_449 (
  .O(douta[29]),
  .I0(mux_o_447),
  .I1(mux_o_448),
  .S0(dff_q_0)
);
MUX2 mux_inst_450 (
  .O(mux_o_450),
  .I0(dpb_inst_16_douta[30]),
  .I1(dpb_inst_17_douta[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_451 (
  .O(mux_o_451),
  .I0(dpb_inst_18_douta[30]),
  .I1(dpb_inst_19_douta[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_452 (
  .O(mux_o_452),
  .I0(dpb_inst_20_douta[30]),
  .I1(dpb_inst_21_douta[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_453 (
  .O(mux_o_453),
  .I0(dpb_inst_22_douta[30]),
  .I1(dpb_inst_23_douta[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_454 (
  .O(mux_o_454),
  .I0(dpb_inst_24_douta[30]),
  .I1(dpb_inst_25_douta[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_455 (
  .O(mux_o_455),
  .I0(dpb_inst_26_douta[30]),
  .I1(dpb_inst_27_douta[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_456 (
  .O(mux_o_456),
  .I0(dpb_inst_28_douta[30]),
  .I1(dpb_inst_29_douta[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_457 (
  .O(mux_o_457),
  .I0(dpb_inst_30_douta[30]),
  .I1(dpb_inst_31_douta[30]),
  .S0(dff_q_3)
);
MUX2 mux_inst_458 (
  .O(mux_o_458),
  .I0(mux_o_450),
  .I1(mux_o_451),
  .S0(dff_q_2)
);
MUX2 mux_inst_459 (
  .O(mux_o_459),
  .I0(mux_o_452),
  .I1(mux_o_453),
  .S0(dff_q_2)
);
MUX2 mux_inst_460 (
  .O(mux_o_460),
  .I0(mux_o_454),
  .I1(mux_o_455),
  .S0(dff_q_2)
);
MUX2 mux_inst_461 (
  .O(mux_o_461),
  .I0(mux_o_456),
  .I1(mux_o_457),
  .S0(dff_q_2)
);
MUX2 mux_inst_462 (
  .O(mux_o_462),
  .I0(mux_o_458),
  .I1(mux_o_459),
  .S0(dff_q_1)
);
MUX2 mux_inst_463 (
  .O(mux_o_463),
  .I0(mux_o_460),
  .I1(mux_o_461),
  .S0(dff_q_1)
);
MUX2 mux_inst_464 (
  .O(douta[30]),
  .I0(mux_o_462),
  .I1(mux_o_463),
  .S0(dff_q_0)
);
MUX2 mux_inst_465 (
  .O(mux_o_465),
  .I0(dpb_inst_16_douta[31]),
  .I1(dpb_inst_17_douta[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_466 (
  .O(mux_o_466),
  .I0(dpb_inst_18_douta[31]),
  .I1(dpb_inst_19_douta[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_467 (
  .O(mux_o_467),
  .I0(dpb_inst_20_douta[31]),
  .I1(dpb_inst_21_douta[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_468 (
  .O(mux_o_468),
  .I0(dpb_inst_22_douta[31]),
  .I1(dpb_inst_23_douta[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_469 (
  .O(mux_o_469),
  .I0(dpb_inst_24_douta[31]),
  .I1(dpb_inst_25_douta[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_470 (
  .O(mux_o_470),
  .I0(dpb_inst_26_douta[31]),
  .I1(dpb_inst_27_douta[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_471 (
  .O(mux_o_471),
  .I0(dpb_inst_28_douta[31]),
  .I1(dpb_inst_29_douta[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_472 (
  .O(mux_o_472),
  .I0(dpb_inst_30_douta[31]),
  .I1(dpb_inst_31_douta[31]),
  .S0(dff_q_3)
);
MUX2 mux_inst_473 (
  .O(mux_o_473),
  .I0(mux_o_465),
  .I1(mux_o_466),
  .S0(dff_q_2)
);
MUX2 mux_inst_474 (
  .O(mux_o_474),
  .I0(mux_o_467),
  .I1(mux_o_468),
  .S0(dff_q_2)
);
MUX2 mux_inst_475 (
  .O(mux_o_475),
  .I0(mux_o_469),
  .I1(mux_o_470),
  .S0(dff_q_2)
);
MUX2 mux_inst_476 (
  .O(mux_o_476),
  .I0(mux_o_471),
  .I1(mux_o_472),
  .S0(dff_q_2)
);
MUX2 mux_inst_477 (
  .O(mux_o_477),
  .I0(mux_o_473),
  .I1(mux_o_474),
  .S0(dff_q_1)
);
MUX2 mux_inst_478 (
  .O(mux_o_478),
  .I0(mux_o_475),
  .I1(mux_o_476),
  .S0(dff_q_1)
);
MUX2 mux_inst_479 (
  .O(douta[31]),
  .I0(mux_o_477),
  .I1(mux_o_478),
  .S0(dff_q_0)
);
MUX2 mux_inst_480 (
  .O(mux_o_480),
  .I0(dpb_inst_0_doutb[0]),
  .I1(dpb_inst_1_doutb[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_481 (
  .O(mux_o_481),
  .I0(dpb_inst_2_doutb[0]),
  .I1(dpb_inst_3_doutb[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_482 (
  .O(mux_o_482),
  .I0(dpb_inst_4_doutb[0]),
  .I1(dpb_inst_5_doutb[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_483 (
  .O(mux_o_483),
  .I0(dpb_inst_6_doutb[0]),
  .I1(dpb_inst_7_doutb[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_484 (
  .O(mux_o_484),
  .I0(dpb_inst_8_doutb[0]),
  .I1(dpb_inst_9_doutb[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_485 (
  .O(mux_o_485),
  .I0(dpb_inst_10_doutb[0]),
  .I1(dpb_inst_11_doutb[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_486 (
  .O(mux_o_486),
  .I0(dpb_inst_12_doutb[0]),
  .I1(dpb_inst_13_doutb[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_487 (
  .O(mux_o_487),
  .I0(dpb_inst_14_doutb[0]),
  .I1(dpb_inst_15_doutb[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_488 (
  .O(mux_o_488),
  .I0(mux_o_480),
  .I1(mux_o_481),
  .S0(dff_q_6)
);
MUX2 mux_inst_489 (
  .O(mux_o_489),
  .I0(mux_o_482),
  .I1(mux_o_483),
  .S0(dff_q_6)
);
MUX2 mux_inst_490 (
  .O(mux_o_490),
  .I0(mux_o_484),
  .I1(mux_o_485),
  .S0(dff_q_6)
);
MUX2 mux_inst_491 (
  .O(mux_o_491),
  .I0(mux_o_486),
  .I1(mux_o_487),
  .S0(dff_q_6)
);
MUX2 mux_inst_492 (
  .O(mux_o_492),
  .I0(mux_o_488),
  .I1(mux_o_489),
  .S0(dff_q_5)
);
MUX2 mux_inst_493 (
  .O(mux_o_493),
  .I0(mux_o_490),
  .I1(mux_o_491),
  .S0(dff_q_5)
);
MUX2 mux_inst_494 (
  .O(doutb[0]),
  .I0(mux_o_492),
  .I1(mux_o_493),
  .S0(dff_q_4)
);
MUX2 mux_inst_495 (
  .O(mux_o_495),
  .I0(dpb_inst_0_doutb[1]),
  .I1(dpb_inst_1_doutb[1]),
  .S0(dff_q_7)
);
MUX2 mux_inst_496 (
  .O(mux_o_496),
  .I0(dpb_inst_2_doutb[1]),
  .I1(dpb_inst_3_doutb[1]),
  .S0(dff_q_7)
);
MUX2 mux_inst_497 (
  .O(mux_o_497),
  .I0(dpb_inst_4_doutb[1]),
  .I1(dpb_inst_5_doutb[1]),
  .S0(dff_q_7)
);
MUX2 mux_inst_498 (
  .O(mux_o_498),
  .I0(dpb_inst_6_doutb[1]),
  .I1(dpb_inst_7_doutb[1]),
  .S0(dff_q_7)
);
MUX2 mux_inst_499 (
  .O(mux_o_499),
  .I0(dpb_inst_8_doutb[1]),
  .I1(dpb_inst_9_doutb[1]),
  .S0(dff_q_7)
);
MUX2 mux_inst_500 (
  .O(mux_o_500),
  .I0(dpb_inst_10_doutb[1]),
  .I1(dpb_inst_11_doutb[1]),
  .S0(dff_q_7)
);
MUX2 mux_inst_501 (
  .O(mux_o_501),
  .I0(dpb_inst_12_doutb[1]),
  .I1(dpb_inst_13_doutb[1]),
  .S0(dff_q_7)
);
MUX2 mux_inst_502 (
  .O(mux_o_502),
  .I0(dpb_inst_14_doutb[1]),
  .I1(dpb_inst_15_doutb[1]),
  .S0(dff_q_7)
);
MUX2 mux_inst_503 (
  .O(mux_o_503),
  .I0(mux_o_495),
  .I1(mux_o_496),
  .S0(dff_q_6)
);
MUX2 mux_inst_504 (
  .O(mux_o_504),
  .I0(mux_o_497),
  .I1(mux_o_498),
  .S0(dff_q_6)
);
MUX2 mux_inst_505 (
  .O(mux_o_505),
  .I0(mux_o_499),
  .I1(mux_o_500),
  .S0(dff_q_6)
);
MUX2 mux_inst_506 (
  .O(mux_o_506),
  .I0(mux_o_501),
  .I1(mux_o_502),
  .S0(dff_q_6)
);
MUX2 mux_inst_507 (
  .O(mux_o_507),
  .I0(mux_o_503),
  .I1(mux_o_504),
  .S0(dff_q_5)
);
MUX2 mux_inst_508 (
  .O(mux_o_508),
  .I0(mux_o_505),
  .I1(mux_o_506),
  .S0(dff_q_5)
);
MUX2 mux_inst_509 (
  .O(doutb[1]),
  .I0(mux_o_507),
  .I1(mux_o_508),
  .S0(dff_q_4)
);
MUX2 mux_inst_510 (
  .O(mux_o_510),
  .I0(dpb_inst_0_doutb[2]),
  .I1(dpb_inst_1_doutb[2]),
  .S0(dff_q_7)
);
MUX2 mux_inst_511 (
  .O(mux_o_511),
  .I0(dpb_inst_2_doutb[2]),
  .I1(dpb_inst_3_doutb[2]),
  .S0(dff_q_7)
);
MUX2 mux_inst_512 (
  .O(mux_o_512),
  .I0(dpb_inst_4_doutb[2]),
  .I1(dpb_inst_5_doutb[2]),
  .S0(dff_q_7)
);
MUX2 mux_inst_513 (
  .O(mux_o_513),
  .I0(dpb_inst_6_doutb[2]),
  .I1(dpb_inst_7_doutb[2]),
  .S0(dff_q_7)
);
MUX2 mux_inst_514 (
  .O(mux_o_514),
  .I0(dpb_inst_8_doutb[2]),
  .I1(dpb_inst_9_doutb[2]),
  .S0(dff_q_7)
);
MUX2 mux_inst_515 (
  .O(mux_o_515),
  .I0(dpb_inst_10_doutb[2]),
  .I1(dpb_inst_11_doutb[2]),
  .S0(dff_q_7)
);
MUX2 mux_inst_516 (
  .O(mux_o_516),
  .I0(dpb_inst_12_doutb[2]),
  .I1(dpb_inst_13_doutb[2]),
  .S0(dff_q_7)
);
MUX2 mux_inst_517 (
  .O(mux_o_517),
  .I0(dpb_inst_14_doutb[2]),
  .I1(dpb_inst_15_doutb[2]),
  .S0(dff_q_7)
);
MUX2 mux_inst_518 (
  .O(mux_o_518),
  .I0(mux_o_510),
  .I1(mux_o_511),
  .S0(dff_q_6)
);
MUX2 mux_inst_519 (
  .O(mux_o_519),
  .I0(mux_o_512),
  .I1(mux_o_513),
  .S0(dff_q_6)
);
MUX2 mux_inst_520 (
  .O(mux_o_520),
  .I0(mux_o_514),
  .I1(mux_o_515),
  .S0(dff_q_6)
);
MUX2 mux_inst_521 (
  .O(mux_o_521),
  .I0(mux_o_516),
  .I1(mux_o_517),
  .S0(dff_q_6)
);
MUX2 mux_inst_522 (
  .O(mux_o_522),
  .I0(mux_o_518),
  .I1(mux_o_519),
  .S0(dff_q_5)
);
MUX2 mux_inst_523 (
  .O(mux_o_523),
  .I0(mux_o_520),
  .I1(mux_o_521),
  .S0(dff_q_5)
);
MUX2 mux_inst_524 (
  .O(doutb[2]),
  .I0(mux_o_522),
  .I1(mux_o_523),
  .S0(dff_q_4)
);
MUX2 mux_inst_525 (
  .O(mux_o_525),
  .I0(dpb_inst_0_doutb[3]),
  .I1(dpb_inst_1_doutb[3]),
  .S0(dff_q_7)
);
MUX2 mux_inst_526 (
  .O(mux_o_526),
  .I0(dpb_inst_2_doutb[3]),
  .I1(dpb_inst_3_doutb[3]),
  .S0(dff_q_7)
);
MUX2 mux_inst_527 (
  .O(mux_o_527),
  .I0(dpb_inst_4_doutb[3]),
  .I1(dpb_inst_5_doutb[3]),
  .S0(dff_q_7)
);
MUX2 mux_inst_528 (
  .O(mux_o_528),
  .I0(dpb_inst_6_doutb[3]),
  .I1(dpb_inst_7_doutb[3]),
  .S0(dff_q_7)
);
MUX2 mux_inst_529 (
  .O(mux_o_529),
  .I0(dpb_inst_8_doutb[3]),
  .I1(dpb_inst_9_doutb[3]),
  .S0(dff_q_7)
);
MUX2 mux_inst_530 (
  .O(mux_o_530),
  .I0(dpb_inst_10_doutb[3]),
  .I1(dpb_inst_11_doutb[3]),
  .S0(dff_q_7)
);
MUX2 mux_inst_531 (
  .O(mux_o_531),
  .I0(dpb_inst_12_doutb[3]),
  .I1(dpb_inst_13_doutb[3]),
  .S0(dff_q_7)
);
MUX2 mux_inst_532 (
  .O(mux_o_532),
  .I0(dpb_inst_14_doutb[3]),
  .I1(dpb_inst_15_doutb[3]),
  .S0(dff_q_7)
);
MUX2 mux_inst_533 (
  .O(mux_o_533),
  .I0(mux_o_525),
  .I1(mux_o_526),
  .S0(dff_q_6)
);
MUX2 mux_inst_534 (
  .O(mux_o_534),
  .I0(mux_o_527),
  .I1(mux_o_528),
  .S0(dff_q_6)
);
MUX2 mux_inst_535 (
  .O(mux_o_535),
  .I0(mux_o_529),
  .I1(mux_o_530),
  .S0(dff_q_6)
);
MUX2 mux_inst_536 (
  .O(mux_o_536),
  .I0(mux_o_531),
  .I1(mux_o_532),
  .S0(dff_q_6)
);
MUX2 mux_inst_537 (
  .O(mux_o_537),
  .I0(mux_o_533),
  .I1(mux_o_534),
  .S0(dff_q_5)
);
MUX2 mux_inst_538 (
  .O(mux_o_538),
  .I0(mux_o_535),
  .I1(mux_o_536),
  .S0(dff_q_5)
);
MUX2 mux_inst_539 (
  .O(doutb[3]),
  .I0(mux_o_537),
  .I1(mux_o_538),
  .S0(dff_q_4)
);
MUX2 mux_inst_540 (
  .O(mux_o_540),
  .I0(dpb_inst_0_doutb[4]),
  .I1(dpb_inst_1_doutb[4]),
  .S0(dff_q_7)
);
MUX2 mux_inst_541 (
  .O(mux_o_541),
  .I0(dpb_inst_2_doutb[4]),
  .I1(dpb_inst_3_doutb[4]),
  .S0(dff_q_7)
);
MUX2 mux_inst_542 (
  .O(mux_o_542),
  .I0(dpb_inst_4_doutb[4]),
  .I1(dpb_inst_5_doutb[4]),
  .S0(dff_q_7)
);
MUX2 mux_inst_543 (
  .O(mux_o_543),
  .I0(dpb_inst_6_doutb[4]),
  .I1(dpb_inst_7_doutb[4]),
  .S0(dff_q_7)
);
MUX2 mux_inst_544 (
  .O(mux_o_544),
  .I0(dpb_inst_8_doutb[4]),
  .I1(dpb_inst_9_doutb[4]),
  .S0(dff_q_7)
);
MUX2 mux_inst_545 (
  .O(mux_o_545),
  .I0(dpb_inst_10_doutb[4]),
  .I1(dpb_inst_11_doutb[4]),
  .S0(dff_q_7)
);
MUX2 mux_inst_546 (
  .O(mux_o_546),
  .I0(dpb_inst_12_doutb[4]),
  .I1(dpb_inst_13_doutb[4]),
  .S0(dff_q_7)
);
MUX2 mux_inst_547 (
  .O(mux_o_547),
  .I0(dpb_inst_14_doutb[4]),
  .I1(dpb_inst_15_doutb[4]),
  .S0(dff_q_7)
);
MUX2 mux_inst_548 (
  .O(mux_o_548),
  .I0(mux_o_540),
  .I1(mux_o_541),
  .S0(dff_q_6)
);
MUX2 mux_inst_549 (
  .O(mux_o_549),
  .I0(mux_o_542),
  .I1(mux_o_543),
  .S0(dff_q_6)
);
MUX2 mux_inst_550 (
  .O(mux_o_550),
  .I0(mux_o_544),
  .I1(mux_o_545),
  .S0(dff_q_6)
);
MUX2 mux_inst_551 (
  .O(mux_o_551),
  .I0(mux_o_546),
  .I1(mux_o_547),
  .S0(dff_q_6)
);
MUX2 mux_inst_552 (
  .O(mux_o_552),
  .I0(mux_o_548),
  .I1(mux_o_549),
  .S0(dff_q_5)
);
MUX2 mux_inst_553 (
  .O(mux_o_553),
  .I0(mux_o_550),
  .I1(mux_o_551),
  .S0(dff_q_5)
);
MUX2 mux_inst_554 (
  .O(doutb[4]),
  .I0(mux_o_552),
  .I1(mux_o_553),
  .S0(dff_q_4)
);
MUX2 mux_inst_555 (
  .O(mux_o_555),
  .I0(dpb_inst_0_doutb[5]),
  .I1(dpb_inst_1_doutb[5]),
  .S0(dff_q_7)
);
MUX2 mux_inst_556 (
  .O(mux_o_556),
  .I0(dpb_inst_2_doutb[5]),
  .I1(dpb_inst_3_doutb[5]),
  .S0(dff_q_7)
);
MUX2 mux_inst_557 (
  .O(mux_o_557),
  .I0(dpb_inst_4_doutb[5]),
  .I1(dpb_inst_5_doutb[5]),
  .S0(dff_q_7)
);
MUX2 mux_inst_558 (
  .O(mux_o_558),
  .I0(dpb_inst_6_doutb[5]),
  .I1(dpb_inst_7_doutb[5]),
  .S0(dff_q_7)
);
MUX2 mux_inst_559 (
  .O(mux_o_559),
  .I0(dpb_inst_8_doutb[5]),
  .I1(dpb_inst_9_doutb[5]),
  .S0(dff_q_7)
);
MUX2 mux_inst_560 (
  .O(mux_o_560),
  .I0(dpb_inst_10_doutb[5]),
  .I1(dpb_inst_11_doutb[5]),
  .S0(dff_q_7)
);
MUX2 mux_inst_561 (
  .O(mux_o_561),
  .I0(dpb_inst_12_doutb[5]),
  .I1(dpb_inst_13_doutb[5]),
  .S0(dff_q_7)
);
MUX2 mux_inst_562 (
  .O(mux_o_562),
  .I0(dpb_inst_14_doutb[5]),
  .I1(dpb_inst_15_doutb[5]),
  .S0(dff_q_7)
);
MUX2 mux_inst_563 (
  .O(mux_o_563),
  .I0(mux_o_555),
  .I1(mux_o_556),
  .S0(dff_q_6)
);
MUX2 mux_inst_564 (
  .O(mux_o_564),
  .I0(mux_o_557),
  .I1(mux_o_558),
  .S0(dff_q_6)
);
MUX2 mux_inst_565 (
  .O(mux_o_565),
  .I0(mux_o_559),
  .I1(mux_o_560),
  .S0(dff_q_6)
);
MUX2 mux_inst_566 (
  .O(mux_o_566),
  .I0(mux_o_561),
  .I1(mux_o_562),
  .S0(dff_q_6)
);
MUX2 mux_inst_567 (
  .O(mux_o_567),
  .I0(mux_o_563),
  .I1(mux_o_564),
  .S0(dff_q_5)
);
MUX2 mux_inst_568 (
  .O(mux_o_568),
  .I0(mux_o_565),
  .I1(mux_o_566),
  .S0(dff_q_5)
);
MUX2 mux_inst_569 (
  .O(doutb[5]),
  .I0(mux_o_567),
  .I1(mux_o_568),
  .S0(dff_q_4)
);
MUX2 mux_inst_570 (
  .O(mux_o_570),
  .I0(dpb_inst_0_doutb[6]),
  .I1(dpb_inst_1_doutb[6]),
  .S0(dff_q_7)
);
MUX2 mux_inst_571 (
  .O(mux_o_571),
  .I0(dpb_inst_2_doutb[6]),
  .I1(dpb_inst_3_doutb[6]),
  .S0(dff_q_7)
);
MUX2 mux_inst_572 (
  .O(mux_o_572),
  .I0(dpb_inst_4_doutb[6]),
  .I1(dpb_inst_5_doutb[6]),
  .S0(dff_q_7)
);
MUX2 mux_inst_573 (
  .O(mux_o_573),
  .I0(dpb_inst_6_doutb[6]),
  .I1(dpb_inst_7_doutb[6]),
  .S0(dff_q_7)
);
MUX2 mux_inst_574 (
  .O(mux_o_574),
  .I0(dpb_inst_8_doutb[6]),
  .I1(dpb_inst_9_doutb[6]),
  .S0(dff_q_7)
);
MUX2 mux_inst_575 (
  .O(mux_o_575),
  .I0(dpb_inst_10_doutb[6]),
  .I1(dpb_inst_11_doutb[6]),
  .S0(dff_q_7)
);
MUX2 mux_inst_576 (
  .O(mux_o_576),
  .I0(dpb_inst_12_doutb[6]),
  .I1(dpb_inst_13_doutb[6]),
  .S0(dff_q_7)
);
MUX2 mux_inst_577 (
  .O(mux_o_577),
  .I0(dpb_inst_14_doutb[6]),
  .I1(dpb_inst_15_doutb[6]),
  .S0(dff_q_7)
);
MUX2 mux_inst_578 (
  .O(mux_o_578),
  .I0(mux_o_570),
  .I1(mux_o_571),
  .S0(dff_q_6)
);
MUX2 mux_inst_579 (
  .O(mux_o_579),
  .I0(mux_o_572),
  .I1(mux_o_573),
  .S0(dff_q_6)
);
MUX2 mux_inst_580 (
  .O(mux_o_580),
  .I0(mux_o_574),
  .I1(mux_o_575),
  .S0(dff_q_6)
);
MUX2 mux_inst_581 (
  .O(mux_o_581),
  .I0(mux_o_576),
  .I1(mux_o_577),
  .S0(dff_q_6)
);
MUX2 mux_inst_582 (
  .O(mux_o_582),
  .I0(mux_o_578),
  .I1(mux_o_579),
  .S0(dff_q_5)
);
MUX2 mux_inst_583 (
  .O(mux_o_583),
  .I0(mux_o_580),
  .I1(mux_o_581),
  .S0(dff_q_5)
);
MUX2 mux_inst_584 (
  .O(doutb[6]),
  .I0(mux_o_582),
  .I1(mux_o_583),
  .S0(dff_q_4)
);
MUX2 mux_inst_585 (
  .O(mux_o_585),
  .I0(dpb_inst_0_doutb[7]),
  .I1(dpb_inst_1_doutb[7]),
  .S0(dff_q_7)
);
MUX2 mux_inst_586 (
  .O(mux_o_586),
  .I0(dpb_inst_2_doutb[7]),
  .I1(dpb_inst_3_doutb[7]),
  .S0(dff_q_7)
);
MUX2 mux_inst_587 (
  .O(mux_o_587),
  .I0(dpb_inst_4_doutb[7]),
  .I1(dpb_inst_5_doutb[7]),
  .S0(dff_q_7)
);
MUX2 mux_inst_588 (
  .O(mux_o_588),
  .I0(dpb_inst_6_doutb[7]),
  .I1(dpb_inst_7_doutb[7]),
  .S0(dff_q_7)
);
MUX2 mux_inst_589 (
  .O(mux_o_589),
  .I0(dpb_inst_8_doutb[7]),
  .I1(dpb_inst_9_doutb[7]),
  .S0(dff_q_7)
);
MUX2 mux_inst_590 (
  .O(mux_o_590),
  .I0(dpb_inst_10_doutb[7]),
  .I1(dpb_inst_11_doutb[7]),
  .S0(dff_q_7)
);
MUX2 mux_inst_591 (
  .O(mux_o_591),
  .I0(dpb_inst_12_doutb[7]),
  .I1(dpb_inst_13_doutb[7]),
  .S0(dff_q_7)
);
MUX2 mux_inst_592 (
  .O(mux_o_592),
  .I0(dpb_inst_14_doutb[7]),
  .I1(dpb_inst_15_doutb[7]),
  .S0(dff_q_7)
);
MUX2 mux_inst_593 (
  .O(mux_o_593),
  .I0(mux_o_585),
  .I1(mux_o_586),
  .S0(dff_q_6)
);
MUX2 mux_inst_594 (
  .O(mux_o_594),
  .I0(mux_o_587),
  .I1(mux_o_588),
  .S0(dff_q_6)
);
MUX2 mux_inst_595 (
  .O(mux_o_595),
  .I0(mux_o_589),
  .I1(mux_o_590),
  .S0(dff_q_6)
);
MUX2 mux_inst_596 (
  .O(mux_o_596),
  .I0(mux_o_591),
  .I1(mux_o_592),
  .S0(dff_q_6)
);
MUX2 mux_inst_597 (
  .O(mux_o_597),
  .I0(mux_o_593),
  .I1(mux_o_594),
  .S0(dff_q_5)
);
MUX2 mux_inst_598 (
  .O(mux_o_598),
  .I0(mux_o_595),
  .I1(mux_o_596),
  .S0(dff_q_5)
);
MUX2 mux_inst_599 (
  .O(doutb[7]),
  .I0(mux_o_597),
  .I1(mux_o_598),
  .S0(dff_q_4)
);
MUX2 mux_inst_600 (
  .O(mux_o_600),
  .I0(dpb_inst_0_doutb[8]),
  .I1(dpb_inst_1_doutb[8]),
  .S0(dff_q_7)
);
MUX2 mux_inst_601 (
  .O(mux_o_601),
  .I0(dpb_inst_2_doutb[8]),
  .I1(dpb_inst_3_doutb[8]),
  .S0(dff_q_7)
);
MUX2 mux_inst_602 (
  .O(mux_o_602),
  .I0(dpb_inst_4_doutb[8]),
  .I1(dpb_inst_5_doutb[8]),
  .S0(dff_q_7)
);
MUX2 mux_inst_603 (
  .O(mux_o_603),
  .I0(dpb_inst_6_doutb[8]),
  .I1(dpb_inst_7_doutb[8]),
  .S0(dff_q_7)
);
MUX2 mux_inst_604 (
  .O(mux_o_604),
  .I0(dpb_inst_8_doutb[8]),
  .I1(dpb_inst_9_doutb[8]),
  .S0(dff_q_7)
);
MUX2 mux_inst_605 (
  .O(mux_o_605),
  .I0(dpb_inst_10_doutb[8]),
  .I1(dpb_inst_11_doutb[8]),
  .S0(dff_q_7)
);
MUX2 mux_inst_606 (
  .O(mux_o_606),
  .I0(dpb_inst_12_doutb[8]),
  .I1(dpb_inst_13_doutb[8]),
  .S0(dff_q_7)
);
MUX2 mux_inst_607 (
  .O(mux_o_607),
  .I0(dpb_inst_14_doutb[8]),
  .I1(dpb_inst_15_doutb[8]),
  .S0(dff_q_7)
);
MUX2 mux_inst_608 (
  .O(mux_o_608),
  .I0(mux_o_600),
  .I1(mux_o_601),
  .S0(dff_q_6)
);
MUX2 mux_inst_609 (
  .O(mux_o_609),
  .I0(mux_o_602),
  .I1(mux_o_603),
  .S0(dff_q_6)
);
MUX2 mux_inst_610 (
  .O(mux_o_610),
  .I0(mux_o_604),
  .I1(mux_o_605),
  .S0(dff_q_6)
);
MUX2 mux_inst_611 (
  .O(mux_o_611),
  .I0(mux_o_606),
  .I1(mux_o_607),
  .S0(dff_q_6)
);
MUX2 mux_inst_612 (
  .O(mux_o_612),
  .I0(mux_o_608),
  .I1(mux_o_609),
  .S0(dff_q_5)
);
MUX2 mux_inst_613 (
  .O(mux_o_613),
  .I0(mux_o_610),
  .I1(mux_o_611),
  .S0(dff_q_5)
);
MUX2 mux_inst_614 (
  .O(doutb[8]),
  .I0(mux_o_612),
  .I1(mux_o_613),
  .S0(dff_q_4)
);
MUX2 mux_inst_615 (
  .O(mux_o_615),
  .I0(dpb_inst_0_doutb[9]),
  .I1(dpb_inst_1_doutb[9]),
  .S0(dff_q_7)
);
MUX2 mux_inst_616 (
  .O(mux_o_616),
  .I0(dpb_inst_2_doutb[9]),
  .I1(dpb_inst_3_doutb[9]),
  .S0(dff_q_7)
);
MUX2 mux_inst_617 (
  .O(mux_o_617),
  .I0(dpb_inst_4_doutb[9]),
  .I1(dpb_inst_5_doutb[9]),
  .S0(dff_q_7)
);
MUX2 mux_inst_618 (
  .O(mux_o_618),
  .I0(dpb_inst_6_doutb[9]),
  .I1(dpb_inst_7_doutb[9]),
  .S0(dff_q_7)
);
MUX2 mux_inst_619 (
  .O(mux_o_619),
  .I0(dpb_inst_8_doutb[9]),
  .I1(dpb_inst_9_doutb[9]),
  .S0(dff_q_7)
);
MUX2 mux_inst_620 (
  .O(mux_o_620),
  .I0(dpb_inst_10_doutb[9]),
  .I1(dpb_inst_11_doutb[9]),
  .S0(dff_q_7)
);
MUX2 mux_inst_621 (
  .O(mux_o_621),
  .I0(dpb_inst_12_doutb[9]),
  .I1(dpb_inst_13_doutb[9]),
  .S0(dff_q_7)
);
MUX2 mux_inst_622 (
  .O(mux_o_622),
  .I0(dpb_inst_14_doutb[9]),
  .I1(dpb_inst_15_doutb[9]),
  .S0(dff_q_7)
);
MUX2 mux_inst_623 (
  .O(mux_o_623),
  .I0(mux_o_615),
  .I1(mux_o_616),
  .S0(dff_q_6)
);
MUX2 mux_inst_624 (
  .O(mux_o_624),
  .I0(mux_o_617),
  .I1(mux_o_618),
  .S0(dff_q_6)
);
MUX2 mux_inst_625 (
  .O(mux_o_625),
  .I0(mux_o_619),
  .I1(mux_o_620),
  .S0(dff_q_6)
);
MUX2 mux_inst_626 (
  .O(mux_o_626),
  .I0(mux_o_621),
  .I1(mux_o_622),
  .S0(dff_q_6)
);
MUX2 mux_inst_627 (
  .O(mux_o_627),
  .I0(mux_o_623),
  .I1(mux_o_624),
  .S0(dff_q_5)
);
MUX2 mux_inst_628 (
  .O(mux_o_628),
  .I0(mux_o_625),
  .I1(mux_o_626),
  .S0(dff_q_5)
);
MUX2 mux_inst_629 (
  .O(doutb[9]),
  .I0(mux_o_627),
  .I1(mux_o_628),
  .S0(dff_q_4)
);
MUX2 mux_inst_630 (
  .O(mux_o_630),
  .I0(dpb_inst_0_doutb[10]),
  .I1(dpb_inst_1_doutb[10]),
  .S0(dff_q_7)
);
MUX2 mux_inst_631 (
  .O(mux_o_631),
  .I0(dpb_inst_2_doutb[10]),
  .I1(dpb_inst_3_doutb[10]),
  .S0(dff_q_7)
);
MUX2 mux_inst_632 (
  .O(mux_o_632),
  .I0(dpb_inst_4_doutb[10]),
  .I1(dpb_inst_5_doutb[10]),
  .S0(dff_q_7)
);
MUX2 mux_inst_633 (
  .O(mux_o_633),
  .I0(dpb_inst_6_doutb[10]),
  .I1(dpb_inst_7_doutb[10]),
  .S0(dff_q_7)
);
MUX2 mux_inst_634 (
  .O(mux_o_634),
  .I0(dpb_inst_8_doutb[10]),
  .I1(dpb_inst_9_doutb[10]),
  .S0(dff_q_7)
);
MUX2 mux_inst_635 (
  .O(mux_o_635),
  .I0(dpb_inst_10_doutb[10]),
  .I1(dpb_inst_11_doutb[10]),
  .S0(dff_q_7)
);
MUX2 mux_inst_636 (
  .O(mux_o_636),
  .I0(dpb_inst_12_doutb[10]),
  .I1(dpb_inst_13_doutb[10]),
  .S0(dff_q_7)
);
MUX2 mux_inst_637 (
  .O(mux_o_637),
  .I0(dpb_inst_14_doutb[10]),
  .I1(dpb_inst_15_doutb[10]),
  .S0(dff_q_7)
);
MUX2 mux_inst_638 (
  .O(mux_o_638),
  .I0(mux_o_630),
  .I1(mux_o_631),
  .S0(dff_q_6)
);
MUX2 mux_inst_639 (
  .O(mux_o_639),
  .I0(mux_o_632),
  .I1(mux_o_633),
  .S0(dff_q_6)
);
MUX2 mux_inst_640 (
  .O(mux_o_640),
  .I0(mux_o_634),
  .I1(mux_o_635),
  .S0(dff_q_6)
);
MUX2 mux_inst_641 (
  .O(mux_o_641),
  .I0(mux_o_636),
  .I1(mux_o_637),
  .S0(dff_q_6)
);
MUX2 mux_inst_642 (
  .O(mux_o_642),
  .I0(mux_o_638),
  .I1(mux_o_639),
  .S0(dff_q_5)
);
MUX2 mux_inst_643 (
  .O(mux_o_643),
  .I0(mux_o_640),
  .I1(mux_o_641),
  .S0(dff_q_5)
);
MUX2 mux_inst_644 (
  .O(doutb[10]),
  .I0(mux_o_642),
  .I1(mux_o_643),
  .S0(dff_q_4)
);
MUX2 mux_inst_645 (
  .O(mux_o_645),
  .I0(dpb_inst_0_doutb[11]),
  .I1(dpb_inst_1_doutb[11]),
  .S0(dff_q_7)
);
MUX2 mux_inst_646 (
  .O(mux_o_646),
  .I0(dpb_inst_2_doutb[11]),
  .I1(dpb_inst_3_doutb[11]),
  .S0(dff_q_7)
);
MUX2 mux_inst_647 (
  .O(mux_o_647),
  .I0(dpb_inst_4_doutb[11]),
  .I1(dpb_inst_5_doutb[11]),
  .S0(dff_q_7)
);
MUX2 mux_inst_648 (
  .O(mux_o_648),
  .I0(dpb_inst_6_doutb[11]),
  .I1(dpb_inst_7_doutb[11]),
  .S0(dff_q_7)
);
MUX2 mux_inst_649 (
  .O(mux_o_649),
  .I0(dpb_inst_8_doutb[11]),
  .I1(dpb_inst_9_doutb[11]),
  .S0(dff_q_7)
);
MUX2 mux_inst_650 (
  .O(mux_o_650),
  .I0(dpb_inst_10_doutb[11]),
  .I1(dpb_inst_11_doutb[11]),
  .S0(dff_q_7)
);
MUX2 mux_inst_651 (
  .O(mux_o_651),
  .I0(dpb_inst_12_doutb[11]),
  .I1(dpb_inst_13_doutb[11]),
  .S0(dff_q_7)
);
MUX2 mux_inst_652 (
  .O(mux_o_652),
  .I0(dpb_inst_14_doutb[11]),
  .I1(dpb_inst_15_doutb[11]),
  .S0(dff_q_7)
);
MUX2 mux_inst_653 (
  .O(mux_o_653),
  .I0(mux_o_645),
  .I1(mux_o_646),
  .S0(dff_q_6)
);
MUX2 mux_inst_654 (
  .O(mux_o_654),
  .I0(mux_o_647),
  .I1(mux_o_648),
  .S0(dff_q_6)
);
MUX2 mux_inst_655 (
  .O(mux_o_655),
  .I0(mux_o_649),
  .I1(mux_o_650),
  .S0(dff_q_6)
);
MUX2 mux_inst_656 (
  .O(mux_o_656),
  .I0(mux_o_651),
  .I1(mux_o_652),
  .S0(dff_q_6)
);
MUX2 mux_inst_657 (
  .O(mux_o_657),
  .I0(mux_o_653),
  .I1(mux_o_654),
  .S0(dff_q_5)
);
MUX2 mux_inst_658 (
  .O(mux_o_658),
  .I0(mux_o_655),
  .I1(mux_o_656),
  .S0(dff_q_5)
);
MUX2 mux_inst_659 (
  .O(doutb[11]),
  .I0(mux_o_657),
  .I1(mux_o_658),
  .S0(dff_q_4)
);
MUX2 mux_inst_660 (
  .O(mux_o_660),
  .I0(dpb_inst_0_doutb[12]),
  .I1(dpb_inst_1_doutb[12]),
  .S0(dff_q_7)
);
MUX2 mux_inst_661 (
  .O(mux_o_661),
  .I0(dpb_inst_2_doutb[12]),
  .I1(dpb_inst_3_doutb[12]),
  .S0(dff_q_7)
);
MUX2 mux_inst_662 (
  .O(mux_o_662),
  .I0(dpb_inst_4_doutb[12]),
  .I1(dpb_inst_5_doutb[12]),
  .S0(dff_q_7)
);
MUX2 mux_inst_663 (
  .O(mux_o_663),
  .I0(dpb_inst_6_doutb[12]),
  .I1(dpb_inst_7_doutb[12]),
  .S0(dff_q_7)
);
MUX2 mux_inst_664 (
  .O(mux_o_664),
  .I0(dpb_inst_8_doutb[12]),
  .I1(dpb_inst_9_doutb[12]),
  .S0(dff_q_7)
);
MUX2 mux_inst_665 (
  .O(mux_o_665),
  .I0(dpb_inst_10_doutb[12]),
  .I1(dpb_inst_11_doutb[12]),
  .S0(dff_q_7)
);
MUX2 mux_inst_666 (
  .O(mux_o_666),
  .I0(dpb_inst_12_doutb[12]),
  .I1(dpb_inst_13_doutb[12]),
  .S0(dff_q_7)
);
MUX2 mux_inst_667 (
  .O(mux_o_667),
  .I0(dpb_inst_14_doutb[12]),
  .I1(dpb_inst_15_doutb[12]),
  .S0(dff_q_7)
);
MUX2 mux_inst_668 (
  .O(mux_o_668),
  .I0(mux_o_660),
  .I1(mux_o_661),
  .S0(dff_q_6)
);
MUX2 mux_inst_669 (
  .O(mux_o_669),
  .I0(mux_o_662),
  .I1(mux_o_663),
  .S0(dff_q_6)
);
MUX2 mux_inst_670 (
  .O(mux_o_670),
  .I0(mux_o_664),
  .I1(mux_o_665),
  .S0(dff_q_6)
);
MUX2 mux_inst_671 (
  .O(mux_o_671),
  .I0(mux_o_666),
  .I1(mux_o_667),
  .S0(dff_q_6)
);
MUX2 mux_inst_672 (
  .O(mux_o_672),
  .I0(mux_o_668),
  .I1(mux_o_669),
  .S0(dff_q_5)
);
MUX2 mux_inst_673 (
  .O(mux_o_673),
  .I0(mux_o_670),
  .I1(mux_o_671),
  .S0(dff_q_5)
);
MUX2 mux_inst_674 (
  .O(doutb[12]),
  .I0(mux_o_672),
  .I1(mux_o_673),
  .S0(dff_q_4)
);
MUX2 mux_inst_675 (
  .O(mux_o_675),
  .I0(dpb_inst_0_doutb[13]),
  .I1(dpb_inst_1_doutb[13]),
  .S0(dff_q_7)
);
MUX2 mux_inst_676 (
  .O(mux_o_676),
  .I0(dpb_inst_2_doutb[13]),
  .I1(dpb_inst_3_doutb[13]),
  .S0(dff_q_7)
);
MUX2 mux_inst_677 (
  .O(mux_o_677),
  .I0(dpb_inst_4_doutb[13]),
  .I1(dpb_inst_5_doutb[13]),
  .S0(dff_q_7)
);
MUX2 mux_inst_678 (
  .O(mux_o_678),
  .I0(dpb_inst_6_doutb[13]),
  .I1(dpb_inst_7_doutb[13]),
  .S0(dff_q_7)
);
MUX2 mux_inst_679 (
  .O(mux_o_679),
  .I0(dpb_inst_8_doutb[13]),
  .I1(dpb_inst_9_doutb[13]),
  .S0(dff_q_7)
);
MUX2 mux_inst_680 (
  .O(mux_o_680),
  .I0(dpb_inst_10_doutb[13]),
  .I1(dpb_inst_11_doutb[13]),
  .S0(dff_q_7)
);
MUX2 mux_inst_681 (
  .O(mux_o_681),
  .I0(dpb_inst_12_doutb[13]),
  .I1(dpb_inst_13_doutb[13]),
  .S0(dff_q_7)
);
MUX2 mux_inst_682 (
  .O(mux_o_682),
  .I0(dpb_inst_14_doutb[13]),
  .I1(dpb_inst_15_doutb[13]),
  .S0(dff_q_7)
);
MUX2 mux_inst_683 (
  .O(mux_o_683),
  .I0(mux_o_675),
  .I1(mux_o_676),
  .S0(dff_q_6)
);
MUX2 mux_inst_684 (
  .O(mux_o_684),
  .I0(mux_o_677),
  .I1(mux_o_678),
  .S0(dff_q_6)
);
MUX2 mux_inst_685 (
  .O(mux_o_685),
  .I0(mux_o_679),
  .I1(mux_o_680),
  .S0(dff_q_6)
);
MUX2 mux_inst_686 (
  .O(mux_o_686),
  .I0(mux_o_681),
  .I1(mux_o_682),
  .S0(dff_q_6)
);
MUX2 mux_inst_687 (
  .O(mux_o_687),
  .I0(mux_o_683),
  .I1(mux_o_684),
  .S0(dff_q_5)
);
MUX2 mux_inst_688 (
  .O(mux_o_688),
  .I0(mux_o_685),
  .I1(mux_o_686),
  .S0(dff_q_5)
);
MUX2 mux_inst_689 (
  .O(doutb[13]),
  .I0(mux_o_687),
  .I1(mux_o_688),
  .S0(dff_q_4)
);
MUX2 mux_inst_690 (
  .O(mux_o_690),
  .I0(dpb_inst_0_doutb[14]),
  .I1(dpb_inst_1_doutb[14]),
  .S0(dff_q_7)
);
MUX2 mux_inst_691 (
  .O(mux_o_691),
  .I0(dpb_inst_2_doutb[14]),
  .I1(dpb_inst_3_doutb[14]),
  .S0(dff_q_7)
);
MUX2 mux_inst_692 (
  .O(mux_o_692),
  .I0(dpb_inst_4_doutb[14]),
  .I1(dpb_inst_5_doutb[14]),
  .S0(dff_q_7)
);
MUX2 mux_inst_693 (
  .O(mux_o_693),
  .I0(dpb_inst_6_doutb[14]),
  .I1(dpb_inst_7_doutb[14]),
  .S0(dff_q_7)
);
MUX2 mux_inst_694 (
  .O(mux_o_694),
  .I0(dpb_inst_8_doutb[14]),
  .I1(dpb_inst_9_doutb[14]),
  .S0(dff_q_7)
);
MUX2 mux_inst_695 (
  .O(mux_o_695),
  .I0(dpb_inst_10_doutb[14]),
  .I1(dpb_inst_11_doutb[14]),
  .S0(dff_q_7)
);
MUX2 mux_inst_696 (
  .O(mux_o_696),
  .I0(dpb_inst_12_doutb[14]),
  .I1(dpb_inst_13_doutb[14]),
  .S0(dff_q_7)
);
MUX2 mux_inst_697 (
  .O(mux_o_697),
  .I0(dpb_inst_14_doutb[14]),
  .I1(dpb_inst_15_doutb[14]),
  .S0(dff_q_7)
);
MUX2 mux_inst_698 (
  .O(mux_o_698),
  .I0(mux_o_690),
  .I1(mux_o_691),
  .S0(dff_q_6)
);
MUX2 mux_inst_699 (
  .O(mux_o_699),
  .I0(mux_o_692),
  .I1(mux_o_693),
  .S0(dff_q_6)
);
MUX2 mux_inst_700 (
  .O(mux_o_700),
  .I0(mux_o_694),
  .I1(mux_o_695),
  .S0(dff_q_6)
);
MUX2 mux_inst_701 (
  .O(mux_o_701),
  .I0(mux_o_696),
  .I1(mux_o_697),
  .S0(dff_q_6)
);
MUX2 mux_inst_702 (
  .O(mux_o_702),
  .I0(mux_o_698),
  .I1(mux_o_699),
  .S0(dff_q_5)
);
MUX2 mux_inst_703 (
  .O(mux_o_703),
  .I0(mux_o_700),
  .I1(mux_o_701),
  .S0(dff_q_5)
);
MUX2 mux_inst_704 (
  .O(doutb[14]),
  .I0(mux_o_702),
  .I1(mux_o_703),
  .S0(dff_q_4)
);
MUX2 mux_inst_705 (
  .O(mux_o_705),
  .I0(dpb_inst_0_doutb[15]),
  .I1(dpb_inst_1_doutb[15]),
  .S0(dff_q_7)
);
MUX2 mux_inst_706 (
  .O(mux_o_706),
  .I0(dpb_inst_2_doutb[15]),
  .I1(dpb_inst_3_doutb[15]),
  .S0(dff_q_7)
);
MUX2 mux_inst_707 (
  .O(mux_o_707),
  .I0(dpb_inst_4_doutb[15]),
  .I1(dpb_inst_5_doutb[15]),
  .S0(dff_q_7)
);
MUX2 mux_inst_708 (
  .O(mux_o_708),
  .I0(dpb_inst_6_doutb[15]),
  .I1(dpb_inst_7_doutb[15]),
  .S0(dff_q_7)
);
MUX2 mux_inst_709 (
  .O(mux_o_709),
  .I0(dpb_inst_8_doutb[15]),
  .I1(dpb_inst_9_doutb[15]),
  .S0(dff_q_7)
);
MUX2 mux_inst_710 (
  .O(mux_o_710),
  .I0(dpb_inst_10_doutb[15]),
  .I1(dpb_inst_11_doutb[15]),
  .S0(dff_q_7)
);
MUX2 mux_inst_711 (
  .O(mux_o_711),
  .I0(dpb_inst_12_doutb[15]),
  .I1(dpb_inst_13_doutb[15]),
  .S0(dff_q_7)
);
MUX2 mux_inst_712 (
  .O(mux_o_712),
  .I0(dpb_inst_14_doutb[15]),
  .I1(dpb_inst_15_doutb[15]),
  .S0(dff_q_7)
);
MUX2 mux_inst_713 (
  .O(mux_o_713),
  .I0(mux_o_705),
  .I1(mux_o_706),
  .S0(dff_q_6)
);
MUX2 mux_inst_714 (
  .O(mux_o_714),
  .I0(mux_o_707),
  .I1(mux_o_708),
  .S0(dff_q_6)
);
MUX2 mux_inst_715 (
  .O(mux_o_715),
  .I0(mux_o_709),
  .I1(mux_o_710),
  .S0(dff_q_6)
);
MUX2 mux_inst_716 (
  .O(mux_o_716),
  .I0(mux_o_711),
  .I1(mux_o_712),
  .S0(dff_q_6)
);
MUX2 mux_inst_717 (
  .O(mux_o_717),
  .I0(mux_o_713),
  .I1(mux_o_714),
  .S0(dff_q_5)
);
MUX2 mux_inst_718 (
  .O(mux_o_718),
  .I0(mux_o_715),
  .I1(mux_o_716),
  .S0(dff_q_5)
);
MUX2 mux_inst_719 (
  .O(doutb[15]),
  .I0(mux_o_717),
  .I1(mux_o_718),
  .S0(dff_q_4)
);
MUX2 mux_inst_720 (
  .O(mux_o_720),
  .I0(dpb_inst_16_doutb[16]),
  .I1(dpb_inst_17_doutb[16]),
  .S0(dff_q_7)
);
MUX2 mux_inst_721 (
  .O(mux_o_721),
  .I0(dpb_inst_18_doutb[16]),
  .I1(dpb_inst_19_doutb[16]),
  .S0(dff_q_7)
);
MUX2 mux_inst_722 (
  .O(mux_o_722),
  .I0(dpb_inst_20_doutb[16]),
  .I1(dpb_inst_21_doutb[16]),
  .S0(dff_q_7)
);
MUX2 mux_inst_723 (
  .O(mux_o_723),
  .I0(dpb_inst_22_doutb[16]),
  .I1(dpb_inst_23_doutb[16]),
  .S0(dff_q_7)
);
MUX2 mux_inst_724 (
  .O(mux_o_724),
  .I0(dpb_inst_24_doutb[16]),
  .I1(dpb_inst_25_doutb[16]),
  .S0(dff_q_7)
);
MUX2 mux_inst_725 (
  .O(mux_o_725),
  .I0(dpb_inst_26_doutb[16]),
  .I1(dpb_inst_27_doutb[16]),
  .S0(dff_q_7)
);
MUX2 mux_inst_726 (
  .O(mux_o_726),
  .I0(dpb_inst_28_doutb[16]),
  .I1(dpb_inst_29_doutb[16]),
  .S0(dff_q_7)
);
MUX2 mux_inst_727 (
  .O(mux_o_727),
  .I0(dpb_inst_30_doutb[16]),
  .I1(dpb_inst_31_doutb[16]),
  .S0(dff_q_7)
);
MUX2 mux_inst_728 (
  .O(mux_o_728),
  .I0(mux_o_720),
  .I1(mux_o_721),
  .S0(dff_q_6)
);
MUX2 mux_inst_729 (
  .O(mux_o_729),
  .I0(mux_o_722),
  .I1(mux_o_723),
  .S0(dff_q_6)
);
MUX2 mux_inst_730 (
  .O(mux_o_730),
  .I0(mux_o_724),
  .I1(mux_o_725),
  .S0(dff_q_6)
);
MUX2 mux_inst_731 (
  .O(mux_o_731),
  .I0(mux_o_726),
  .I1(mux_o_727),
  .S0(dff_q_6)
);
MUX2 mux_inst_732 (
  .O(mux_o_732),
  .I0(mux_o_728),
  .I1(mux_o_729),
  .S0(dff_q_5)
);
MUX2 mux_inst_733 (
  .O(mux_o_733),
  .I0(mux_o_730),
  .I1(mux_o_731),
  .S0(dff_q_5)
);
MUX2 mux_inst_734 (
  .O(doutb[16]),
  .I0(mux_o_732),
  .I1(mux_o_733),
  .S0(dff_q_4)
);
MUX2 mux_inst_735 (
  .O(mux_o_735),
  .I0(dpb_inst_16_doutb[17]),
  .I1(dpb_inst_17_doutb[17]),
  .S0(dff_q_7)
);
MUX2 mux_inst_736 (
  .O(mux_o_736),
  .I0(dpb_inst_18_doutb[17]),
  .I1(dpb_inst_19_doutb[17]),
  .S0(dff_q_7)
);
MUX2 mux_inst_737 (
  .O(mux_o_737),
  .I0(dpb_inst_20_doutb[17]),
  .I1(dpb_inst_21_doutb[17]),
  .S0(dff_q_7)
);
MUX2 mux_inst_738 (
  .O(mux_o_738),
  .I0(dpb_inst_22_doutb[17]),
  .I1(dpb_inst_23_doutb[17]),
  .S0(dff_q_7)
);
MUX2 mux_inst_739 (
  .O(mux_o_739),
  .I0(dpb_inst_24_doutb[17]),
  .I1(dpb_inst_25_doutb[17]),
  .S0(dff_q_7)
);
MUX2 mux_inst_740 (
  .O(mux_o_740),
  .I0(dpb_inst_26_doutb[17]),
  .I1(dpb_inst_27_doutb[17]),
  .S0(dff_q_7)
);
MUX2 mux_inst_741 (
  .O(mux_o_741),
  .I0(dpb_inst_28_doutb[17]),
  .I1(dpb_inst_29_doutb[17]),
  .S0(dff_q_7)
);
MUX2 mux_inst_742 (
  .O(mux_o_742),
  .I0(dpb_inst_30_doutb[17]),
  .I1(dpb_inst_31_doutb[17]),
  .S0(dff_q_7)
);
MUX2 mux_inst_743 (
  .O(mux_o_743),
  .I0(mux_o_735),
  .I1(mux_o_736),
  .S0(dff_q_6)
);
MUX2 mux_inst_744 (
  .O(mux_o_744),
  .I0(mux_o_737),
  .I1(mux_o_738),
  .S0(dff_q_6)
);
MUX2 mux_inst_745 (
  .O(mux_o_745),
  .I0(mux_o_739),
  .I1(mux_o_740),
  .S0(dff_q_6)
);
MUX2 mux_inst_746 (
  .O(mux_o_746),
  .I0(mux_o_741),
  .I1(mux_o_742),
  .S0(dff_q_6)
);
MUX2 mux_inst_747 (
  .O(mux_o_747),
  .I0(mux_o_743),
  .I1(mux_o_744),
  .S0(dff_q_5)
);
MUX2 mux_inst_748 (
  .O(mux_o_748),
  .I0(mux_o_745),
  .I1(mux_o_746),
  .S0(dff_q_5)
);
MUX2 mux_inst_749 (
  .O(doutb[17]),
  .I0(mux_o_747),
  .I1(mux_o_748),
  .S0(dff_q_4)
);
MUX2 mux_inst_750 (
  .O(mux_o_750),
  .I0(dpb_inst_16_doutb[18]),
  .I1(dpb_inst_17_doutb[18]),
  .S0(dff_q_7)
);
MUX2 mux_inst_751 (
  .O(mux_o_751),
  .I0(dpb_inst_18_doutb[18]),
  .I1(dpb_inst_19_doutb[18]),
  .S0(dff_q_7)
);
MUX2 mux_inst_752 (
  .O(mux_o_752),
  .I0(dpb_inst_20_doutb[18]),
  .I1(dpb_inst_21_doutb[18]),
  .S0(dff_q_7)
);
MUX2 mux_inst_753 (
  .O(mux_o_753),
  .I0(dpb_inst_22_doutb[18]),
  .I1(dpb_inst_23_doutb[18]),
  .S0(dff_q_7)
);
MUX2 mux_inst_754 (
  .O(mux_o_754),
  .I0(dpb_inst_24_doutb[18]),
  .I1(dpb_inst_25_doutb[18]),
  .S0(dff_q_7)
);
MUX2 mux_inst_755 (
  .O(mux_o_755),
  .I0(dpb_inst_26_doutb[18]),
  .I1(dpb_inst_27_doutb[18]),
  .S0(dff_q_7)
);
MUX2 mux_inst_756 (
  .O(mux_o_756),
  .I0(dpb_inst_28_doutb[18]),
  .I1(dpb_inst_29_doutb[18]),
  .S0(dff_q_7)
);
MUX2 mux_inst_757 (
  .O(mux_o_757),
  .I0(dpb_inst_30_doutb[18]),
  .I1(dpb_inst_31_doutb[18]),
  .S0(dff_q_7)
);
MUX2 mux_inst_758 (
  .O(mux_o_758),
  .I0(mux_o_750),
  .I1(mux_o_751),
  .S0(dff_q_6)
);
MUX2 mux_inst_759 (
  .O(mux_o_759),
  .I0(mux_o_752),
  .I1(mux_o_753),
  .S0(dff_q_6)
);
MUX2 mux_inst_760 (
  .O(mux_o_760),
  .I0(mux_o_754),
  .I1(mux_o_755),
  .S0(dff_q_6)
);
MUX2 mux_inst_761 (
  .O(mux_o_761),
  .I0(mux_o_756),
  .I1(mux_o_757),
  .S0(dff_q_6)
);
MUX2 mux_inst_762 (
  .O(mux_o_762),
  .I0(mux_o_758),
  .I1(mux_o_759),
  .S0(dff_q_5)
);
MUX2 mux_inst_763 (
  .O(mux_o_763),
  .I0(mux_o_760),
  .I1(mux_o_761),
  .S0(dff_q_5)
);
MUX2 mux_inst_764 (
  .O(doutb[18]),
  .I0(mux_o_762),
  .I1(mux_o_763),
  .S0(dff_q_4)
);
MUX2 mux_inst_765 (
  .O(mux_o_765),
  .I0(dpb_inst_16_doutb[19]),
  .I1(dpb_inst_17_doutb[19]),
  .S0(dff_q_7)
);
MUX2 mux_inst_766 (
  .O(mux_o_766),
  .I0(dpb_inst_18_doutb[19]),
  .I1(dpb_inst_19_doutb[19]),
  .S0(dff_q_7)
);
MUX2 mux_inst_767 (
  .O(mux_o_767),
  .I0(dpb_inst_20_doutb[19]),
  .I1(dpb_inst_21_doutb[19]),
  .S0(dff_q_7)
);
MUX2 mux_inst_768 (
  .O(mux_o_768),
  .I0(dpb_inst_22_doutb[19]),
  .I1(dpb_inst_23_doutb[19]),
  .S0(dff_q_7)
);
MUX2 mux_inst_769 (
  .O(mux_o_769),
  .I0(dpb_inst_24_doutb[19]),
  .I1(dpb_inst_25_doutb[19]),
  .S0(dff_q_7)
);
MUX2 mux_inst_770 (
  .O(mux_o_770),
  .I0(dpb_inst_26_doutb[19]),
  .I1(dpb_inst_27_doutb[19]),
  .S0(dff_q_7)
);
MUX2 mux_inst_771 (
  .O(mux_o_771),
  .I0(dpb_inst_28_doutb[19]),
  .I1(dpb_inst_29_doutb[19]),
  .S0(dff_q_7)
);
MUX2 mux_inst_772 (
  .O(mux_o_772),
  .I0(dpb_inst_30_doutb[19]),
  .I1(dpb_inst_31_doutb[19]),
  .S0(dff_q_7)
);
MUX2 mux_inst_773 (
  .O(mux_o_773),
  .I0(mux_o_765),
  .I1(mux_o_766),
  .S0(dff_q_6)
);
MUX2 mux_inst_774 (
  .O(mux_o_774),
  .I0(mux_o_767),
  .I1(mux_o_768),
  .S0(dff_q_6)
);
MUX2 mux_inst_775 (
  .O(mux_o_775),
  .I0(mux_o_769),
  .I1(mux_o_770),
  .S0(dff_q_6)
);
MUX2 mux_inst_776 (
  .O(mux_o_776),
  .I0(mux_o_771),
  .I1(mux_o_772),
  .S0(dff_q_6)
);
MUX2 mux_inst_777 (
  .O(mux_o_777),
  .I0(mux_o_773),
  .I1(mux_o_774),
  .S0(dff_q_5)
);
MUX2 mux_inst_778 (
  .O(mux_o_778),
  .I0(mux_o_775),
  .I1(mux_o_776),
  .S0(dff_q_5)
);
MUX2 mux_inst_779 (
  .O(doutb[19]),
  .I0(mux_o_777),
  .I1(mux_o_778),
  .S0(dff_q_4)
);
MUX2 mux_inst_780 (
  .O(mux_o_780),
  .I0(dpb_inst_16_doutb[20]),
  .I1(dpb_inst_17_doutb[20]),
  .S0(dff_q_7)
);
MUX2 mux_inst_781 (
  .O(mux_o_781),
  .I0(dpb_inst_18_doutb[20]),
  .I1(dpb_inst_19_doutb[20]),
  .S0(dff_q_7)
);
MUX2 mux_inst_782 (
  .O(mux_o_782),
  .I0(dpb_inst_20_doutb[20]),
  .I1(dpb_inst_21_doutb[20]),
  .S0(dff_q_7)
);
MUX2 mux_inst_783 (
  .O(mux_o_783),
  .I0(dpb_inst_22_doutb[20]),
  .I1(dpb_inst_23_doutb[20]),
  .S0(dff_q_7)
);
MUX2 mux_inst_784 (
  .O(mux_o_784),
  .I0(dpb_inst_24_doutb[20]),
  .I1(dpb_inst_25_doutb[20]),
  .S0(dff_q_7)
);
MUX2 mux_inst_785 (
  .O(mux_o_785),
  .I0(dpb_inst_26_doutb[20]),
  .I1(dpb_inst_27_doutb[20]),
  .S0(dff_q_7)
);
MUX2 mux_inst_786 (
  .O(mux_o_786),
  .I0(dpb_inst_28_doutb[20]),
  .I1(dpb_inst_29_doutb[20]),
  .S0(dff_q_7)
);
MUX2 mux_inst_787 (
  .O(mux_o_787),
  .I0(dpb_inst_30_doutb[20]),
  .I1(dpb_inst_31_doutb[20]),
  .S0(dff_q_7)
);
MUX2 mux_inst_788 (
  .O(mux_o_788),
  .I0(mux_o_780),
  .I1(mux_o_781),
  .S0(dff_q_6)
);
MUX2 mux_inst_789 (
  .O(mux_o_789),
  .I0(mux_o_782),
  .I1(mux_o_783),
  .S0(dff_q_6)
);
MUX2 mux_inst_790 (
  .O(mux_o_790),
  .I0(mux_o_784),
  .I1(mux_o_785),
  .S0(dff_q_6)
);
MUX2 mux_inst_791 (
  .O(mux_o_791),
  .I0(mux_o_786),
  .I1(mux_o_787),
  .S0(dff_q_6)
);
MUX2 mux_inst_792 (
  .O(mux_o_792),
  .I0(mux_o_788),
  .I1(mux_o_789),
  .S0(dff_q_5)
);
MUX2 mux_inst_793 (
  .O(mux_o_793),
  .I0(mux_o_790),
  .I1(mux_o_791),
  .S0(dff_q_5)
);
MUX2 mux_inst_794 (
  .O(doutb[20]),
  .I0(mux_o_792),
  .I1(mux_o_793),
  .S0(dff_q_4)
);
MUX2 mux_inst_795 (
  .O(mux_o_795),
  .I0(dpb_inst_16_doutb[21]),
  .I1(dpb_inst_17_doutb[21]),
  .S0(dff_q_7)
);
MUX2 mux_inst_796 (
  .O(mux_o_796),
  .I0(dpb_inst_18_doutb[21]),
  .I1(dpb_inst_19_doutb[21]),
  .S0(dff_q_7)
);
MUX2 mux_inst_797 (
  .O(mux_o_797),
  .I0(dpb_inst_20_doutb[21]),
  .I1(dpb_inst_21_doutb[21]),
  .S0(dff_q_7)
);
MUX2 mux_inst_798 (
  .O(mux_o_798),
  .I0(dpb_inst_22_doutb[21]),
  .I1(dpb_inst_23_doutb[21]),
  .S0(dff_q_7)
);
MUX2 mux_inst_799 (
  .O(mux_o_799),
  .I0(dpb_inst_24_doutb[21]),
  .I1(dpb_inst_25_doutb[21]),
  .S0(dff_q_7)
);
MUX2 mux_inst_800 (
  .O(mux_o_800),
  .I0(dpb_inst_26_doutb[21]),
  .I1(dpb_inst_27_doutb[21]),
  .S0(dff_q_7)
);
MUX2 mux_inst_801 (
  .O(mux_o_801),
  .I0(dpb_inst_28_doutb[21]),
  .I1(dpb_inst_29_doutb[21]),
  .S0(dff_q_7)
);
MUX2 mux_inst_802 (
  .O(mux_o_802),
  .I0(dpb_inst_30_doutb[21]),
  .I1(dpb_inst_31_doutb[21]),
  .S0(dff_q_7)
);
MUX2 mux_inst_803 (
  .O(mux_o_803),
  .I0(mux_o_795),
  .I1(mux_o_796),
  .S0(dff_q_6)
);
MUX2 mux_inst_804 (
  .O(mux_o_804),
  .I0(mux_o_797),
  .I1(mux_o_798),
  .S0(dff_q_6)
);
MUX2 mux_inst_805 (
  .O(mux_o_805),
  .I0(mux_o_799),
  .I1(mux_o_800),
  .S0(dff_q_6)
);
MUX2 mux_inst_806 (
  .O(mux_o_806),
  .I0(mux_o_801),
  .I1(mux_o_802),
  .S0(dff_q_6)
);
MUX2 mux_inst_807 (
  .O(mux_o_807),
  .I0(mux_o_803),
  .I1(mux_o_804),
  .S0(dff_q_5)
);
MUX2 mux_inst_808 (
  .O(mux_o_808),
  .I0(mux_o_805),
  .I1(mux_o_806),
  .S0(dff_q_5)
);
MUX2 mux_inst_809 (
  .O(doutb[21]),
  .I0(mux_o_807),
  .I1(mux_o_808),
  .S0(dff_q_4)
);
MUX2 mux_inst_810 (
  .O(mux_o_810),
  .I0(dpb_inst_16_doutb[22]),
  .I1(dpb_inst_17_doutb[22]),
  .S0(dff_q_7)
);
MUX2 mux_inst_811 (
  .O(mux_o_811),
  .I0(dpb_inst_18_doutb[22]),
  .I1(dpb_inst_19_doutb[22]),
  .S0(dff_q_7)
);
MUX2 mux_inst_812 (
  .O(mux_o_812),
  .I0(dpb_inst_20_doutb[22]),
  .I1(dpb_inst_21_doutb[22]),
  .S0(dff_q_7)
);
MUX2 mux_inst_813 (
  .O(mux_o_813),
  .I0(dpb_inst_22_doutb[22]),
  .I1(dpb_inst_23_doutb[22]),
  .S0(dff_q_7)
);
MUX2 mux_inst_814 (
  .O(mux_o_814),
  .I0(dpb_inst_24_doutb[22]),
  .I1(dpb_inst_25_doutb[22]),
  .S0(dff_q_7)
);
MUX2 mux_inst_815 (
  .O(mux_o_815),
  .I0(dpb_inst_26_doutb[22]),
  .I1(dpb_inst_27_doutb[22]),
  .S0(dff_q_7)
);
MUX2 mux_inst_816 (
  .O(mux_o_816),
  .I0(dpb_inst_28_doutb[22]),
  .I1(dpb_inst_29_doutb[22]),
  .S0(dff_q_7)
);
MUX2 mux_inst_817 (
  .O(mux_o_817),
  .I0(dpb_inst_30_doutb[22]),
  .I1(dpb_inst_31_doutb[22]),
  .S0(dff_q_7)
);
MUX2 mux_inst_818 (
  .O(mux_o_818),
  .I0(mux_o_810),
  .I1(mux_o_811),
  .S0(dff_q_6)
);
MUX2 mux_inst_819 (
  .O(mux_o_819),
  .I0(mux_o_812),
  .I1(mux_o_813),
  .S0(dff_q_6)
);
MUX2 mux_inst_820 (
  .O(mux_o_820),
  .I0(mux_o_814),
  .I1(mux_o_815),
  .S0(dff_q_6)
);
MUX2 mux_inst_821 (
  .O(mux_o_821),
  .I0(mux_o_816),
  .I1(mux_o_817),
  .S0(dff_q_6)
);
MUX2 mux_inst_822 (
  .O(mux_o_822),
  .I0(mux_o_818),
  .I1(mux_o_819),
  .S0(dff_q_5)
);
MUX2 mux_inst_823 (
  .O(mux_o_823),
  .I0(mux_o_820),
  .I1(mux_o_821),
  .S0(dff_q_5)
);
MUX2 mux_inst_824 (
  .O(doutb[22]),
  .I0(mux_o_822),
  .I1(mux_o_823),
  .S0(dff_q_4)
);
MUX2 mux_inst_825 (
  .O(mux_o_825),
  .I0(dpb_inst_16_doutb[23]),
  .I1(dpb_inst_17_doutb[23]),
  .S0(dff_q_7)
);
MUX2 mux_inst_826 (
  .O(mux_o_826),
  .I0(dpb_inst_18_doutb[23]),
  .I1(dpb_inst_19_doutb[23]),
  .S0(dff_q_7)
);
MUX2 mux_inst_827 (
  .O(mux_o_827),
  .I0(dpb_inst_20_doutb[23]),
  .I1(dpb_inst_21_doutb[23]),
  .S0(dff_q_7)
);
MUX2 mux_inst_828 (
  .O(mux_o_828),
  .I0(dpb_inst_22_doutb[23]),
  .I1(dpb_inst_23_doutb[23]),
  .S0(dff_q_7)
);
MUX2 mux_inst_829 (
  .O(mux_o_829),
  .I0(dpb_inst_24_doutb[23]),
  .I1(dpb_inst_25_doutb[23]),
  .S0(dff_q_7)
);
MUX2 mux_inst_830 (
  .O(mux_o_830),
  .I0(dpb_inst_26_doutb[23]),
  .I1(dpb_inst_27_doutb[23]),
  .S0(dff_q_7)
);
MUX2 mux_inst_831 (
  .O(mux_o_831),
  .I0(dpb_inst_28_doutb[23]),
  .I1(dpb_inst_29_doutb[23]),
  .S0(dff_q_7)
);
MUX2 mux_inst_832 (
  .O(mux_o_832),
  .I0(dpb_inst_30_doutb[23]),
  .I1(dpb_inst_31_doutb[23]),
  .S0(dff_q_7)
);
MUX2 mux_inst_833 (
  .O(mux_o_833),
  .I0(mux_o_825),
  .I1(mux_o_826),
  .S0(dff_q_6)
);
MUX2 mux_inst_834 (
  .O(mux_o_834),
  .I0(mux_o_827),
  .I1(mux_o_828),
  .S0(dff_q_6)
);
MUX2 mux_inst_835 (
  .O(mux_o_835),
  .I0(mux_o_829),
  .I1(mux_o_830),
  .S0(dff_q_6)
);
MUX2 mux_inst_836 (
  .O(mux_o_836),
  .I0(mux_o_831),
  .I1(mux_o_832),
  .S0(dff_q_6)
);
MUX2 mux_inst_837 (
  .O(mux_o_837),
  .I0(mux_o_833),
  .I1(mux_o_834),
  .S0(dff_q_5)
);
MUX2 mux_inst_838 (
  .O(mux_o_838),
  .I0(mux_o_835),
  .I1(mux_o_836),
  .S0(dff_q_5)
);
MUX2 mux_inst_839 (
  .O(doutb[23]),
  .I0(mux_o_837),
  .I1(mux_o_838),
  .S0(dff_q_4)
);
MUX2 mux_inst_840 (
  .O(mux_o_840),
  .I0(dpb_inst_16_doutb[24]),
  .I1(dpb_inst_17_doutb[24]),
  .S0(dff_q_7)
);
MUX2 mux_inst_841 (
  .O(mux_o_841),
  .I0(dpb_inst_18_doutb[24]),
  .I1(dpb_inst_19_doutb[24]),
  .S0(dff_q_7)
);
MUX2 mux_inst_842 (
  .O(mux_o_842),
  .I0(dpb_inst_20_doutb[24]),
  .I1(dpb_inst_21_doutb[24]),
  .S0(dff_q_7)
);
MUX2 mux_inst_843 (
  .O(mux_o_843),
  .I0(dpb_inst_22_doutb[24]),
  .I1(dpb_inst_23_doutb[24]),
  .S0(dff_q_7)
);
MUX2 mux_inst_844 (
  .O(mux_o_844),
  .I0(dpb_inst_24_doutb[24]),
  .I1(dpb_inst_25_doutb[24]),
  .S0(dff_q_7)
);
MUX2 mux_inst_845 (
  .O(mux_o_845),
  .I0(dpb_inst_26_doutb[24]),
  .I1(dpb_inst_27_doutb[24]),
  .S0(dff_q_7)
);
MUX2 mux_inst_846 (
  .O(mux_o_846),
  .I0(dpb_inst_28_doutb[24]),
  .I1(dpb_inst_29_doutb[24]),
  .S0(dff_q_7)
);
MUX2 mux_inst_847 (
  .O(mux_o_847),
  .I0(dpb_inst_30_doutb[24]),
  .I1(dpb_inst_31_doutb[24]),
  .S0(dff_q_7)
);
MUX2 mux_inst_848 (
  .O(mux_o_848),
  .I0(mux_o_840),
  .I1(mux_o_841),
  .S0(dff_q_6)
);
MUX2 mux_inst_849 (
  .O(mux_o_849),
  .I0(mux_o_842),
  .I1(mux_o_843),
  .S0(dff_q_6)
);
MUX2 mux_inst_850 (
  .O(mux_o_850),
  .I0(mux_o_844),
  .I1(mux_o_845),
  .S0(dff_q_6)
);
MUX2 mux_inst_851 (
  .O(mux_o_851),
  .I0(mux_o_846),
  .I1(mux_o_847),
  .S0(dff_q_6)
);
MUX2 mux_inst_852 (
  .O(mux_o_852),
  .I0(mux_o_848),
  .I1(mux_o_849),
  .S0(dff_q_5)
);
MUX2 mux_inst_853 (
  .O(mux_o_853),
  .I0(mux_o_850),
  .I1(mux_o_851),
  .S0(dff_q_5)
);
MUX2 mux_inst_854 (
  .O(doutb[24]),
  .I0(mux_o_852),
  .I1(mux_o_853),
  .S0(dff_q_4)
);
MUX2 mux_inst_855 (
  .O(mux_o_855),
  .I0(dpb_inst_16_doutb[25]),
  .I1(dpb_inst_17_doutb[25]),
  .S0(dff_q_7)
);
MUX2 mux_inst_856 (
  .O(mux_o_856),
  .I0(dpb_inst_18_doutb[25]),
  .I1(dpb_inst_19_doutb[25]),
  .S0(dff_q_7)
);
MUX2 mux_inst_857 (
  .O(mux_o_857),
  .I0(dpb_inst_20_doutb[25]),
  .I1(dpb_inst_21_doutb[25]),
  .S0(dff_q_7)
);
MUX2 mux_inst_858 (
  .O(mux_o_858),
  .I0(dpb_inst_22_doutb[25]),
  .I1(dpb_inst_23_doutb[25]),
  .S0(dff_q_7)
);
MUX2 mux_inst_859 (
  .O(mux_o_859),
  .I0(dpb_inst_24_doutb[25]),
  .I1(dpb_inst_25_doutb[25]),
  .S0(dff_q_7)
);
MUX2 mux_inst_860 (
  .O(mux_o_860),
  .I0(dpb_inst_26_doutb[25]),
  .I1(dpb_inst_27_doutb[25]),
  .S0(dff_q_7)
);
MUX2 mux_inst_861 (
  .O(mux_o_861),
  .I0(dpb_inst_28_doutb[25]),
  .I1(dpb_inst_29_doutb[25]),
  .S0(dff_q_7)
);
MUX2 mux_inst_862 (
  .O(mux_o_862),
  .I0(dpb_inst_30_doutb[25]),
  .I1(dpb_inst_31_doutb[25]),
  .S0(dff_q_7)
);
MUX2 mux_inst_863 (
  .O(mux_o_863),
  .I0(mux_o_855),
  .I1(mux_o_856),
  .S0(dff_q_6)
);
MUX2 mux_inst_864 (
  .O(mux_o_864),
  .I0(mux_o_857),
  .I1(mux_o_858),
  .S0(dff_q_6)
);
MUX2 mux_inst_865 (
  .O(mux_o_865),
  .I0(mux_o_859),
  .I1(mux_o_860),
  .S0(dff_q_6)
);
MUX2 mux_inst_866 (
  .O(mux_o_866),
  .I0(mux_o_861),
  .I1(mux_o_862),
  .S0(dff_q_6)
);
MUX2 mux_inst_867 (
  .O(mux_o_867),
  .I0(mux_o_863),
  .I1(mux_o_864),
  .S0(dff_q_5)
);
MUX2 mux_inst_868 (
  .O(mux_o_868),
  .I0(mux_o_865),
  .I1(mux_o_866),
  .S0(dff_q_5)
);
MUX2 mux_inst_869 (
  .O(doutb[25]),
  .I0(mux_o_867),
  .I1(mux_o_868),
  .S0(dff_q_4)
);
MUX2 mux_inst_870 (
  .O(mux_o_870),
  .I0(dpb_inst_16_doutb[26]),
  .I1(dpb_inst_17_doutb[26]),
  .S0(dff_q_7)
);
MUX2 mux_inst_871 (
  .O(mux_o_871),
  .I0(dpb_inst_18_doutb[26]),
  .I1(dpb_inst_19_doutb[26]),
  .S0(dff_q_7)
);
MUX2 mux_inst_872 (
  .O(mux_o_872),
  .I0(dpb_inst_20_doutb[26]),
  .I1(dpb_inst_21_doutb[26]),
  .S0(dff_q_7)
);
MUX2 mux_inst_873 (
  .O(mux_o_873),
  .I0(dpb_inst_22_doutb[26]),
  .I1(dpb_inst_23_doutb[26]),
  .S0(dff_q_7)
);
MUX2 mux_inst_874 (
  .O(mux_o_874),
  .I0(dpb_inst_24_doutb[26]),
  .I1(dpb_inst_25_doutb[26]),
  .S0(dff_q_7)
);
MUX2 mux_inst_875 (
  .O(mux_o_875),
  .I0(dpb_inst_26_doutb[26]),
  .I1(dpb_inst_27_doutb[26]),
  .S0(dff_q_7)
);
MUX2 mux_inst_876 (
  .O(mux_o_876),
  .I0(dpb_inst_28_doutb[26]),
  .I1(dpb_inst_29_doutb[26]),
  .S0(dff_q_7)
);
MUX2 mux_inst_877 (
  .O(mux_o_877),
  .I0(dpb_inst_30_doutb[26]),
  .I1(dpb_inst_31_doutb[26]),
  .S0(dff_q_7)
);
MUX2 mux_inst_878 (
  .O(mux_o_878),
  .I0(mux_o_870),
  .I1(mux_o_871),
  .S0(dff_q_6)
);
MUX2 mux_inst_879 (
  .O(mux_o_879),
  .I0(mux_o_872),
  .I1(mux_o_873),
  .S0(dff_q_6)
);
MUX2 mux_inst_880 (
  .O(mux_o_880),
  .I0(mux_o_874),
  .I1(mux_o_875),
  .S0(dff_q_6)
);
MUX2 mux_inst_881 (
  .O(mux_o_881),
  .I0(mux_o_876),
  .I1(mux_o_877),
  .S0(dff_q_6)
);
MUX2 mux_inst_882 (
  .O(mux_o_882),
  .I0(mux_o_878),
  .I1(mux_o_879),
  .S0(dff_q_5)
);
MUX2 mux_inst_883 (
  .O(mux_o_883),
  .I0(mux_o_880),
  .I1(mux_o_881),
  .S0(dff_q_5)
);
MUX2 mux_inst_884 (
  .O(doutb[26]),
  .I0(mux_o_882),
  .I1(mux_o_883),
  .S0(dff_q_4)
);
MUX2 mux_inst_885 (
  .O(mux_o_885),
  .I0(dpb_inst_16_doutb[27]),
  .I1(dpb_inst_17_doutb[27]),
  .S0(dff_q_7)
);
MUX2 mux_inst_886 (
  .O(mux_o_886),
  .I0(dpb_inst_18_doutb[27]),
  .I1(dpb_inst_19_doutb[27]),
  .S0(dff_q_7)
);
MUX2 mux_inst_887 (
  .O(mux_o_887),
  .I0(dpb_inst_20_doutb[27]),
  .I1(dpb_inst_21_doutb[27]),
  .S0(dff_q_7)
);
MUX2 mux_inst_888 (
  .O(mux_o_888),
  .I0(dpb_inst_22_doutb[27]),
  .I1(dpb_inst_23_doutb[27]),
  .S0(dff_q_7)
);
MUX2 mux_inst_889 (
  .O(mux_o_889),
  .I0(dpb_inst_24_doutb[27]),
  .I1(dpb_inst_25_doutb[27]),
  .S0(dff_q_7)
);
MUX2 mux_inst_890 (
  .O(mux_o_890),
  .I0(dpb_inst_26_doutb[27]),
  .I1(dpb_inst_27_doutb[27]),
  .S0(dff_q_7)
);
MUX2 mux_inst_891 (
  .O(mux_o_891),
  .I0(dpb_inst_28_doutb[27]),
  .I1(dpb_inst_29_doutb[27]),
  .S0(dff_q_7)
);
MUX2 mux_inst_892 (
  .O(mux_o_892),
  .I0(dpb_inst_30_doutb[27]),
  .I1(dpb_inst_31_doutb[27]),
  .S0(dff_q_7)
);
MUX2 mux_inst_893 (
  .O(mux_o_893),
  .I0(mux_o_885),
  .I1(mux_o_886),
  .S0(dff_q_6)
);
MUX2 mux_inst_894 (
  .O(mux_o_894),
  .I0(mux_o_887),
  .I1(mux_o_888),
  .S0(dff_q_6)
);
MUX2 mux_inst_895 (
  .O(mux_o_895),
  .I0(mux_o_889),
  .I1(mux_o_890),
  .S0(dff_q_6)
);
MUX2 mux_inst_896 (
  .O(mux_o_896),
  .I0(mux_o_891),
  .I1(mux_o_892),
  .S0(dff_q_6)
);
MUX2 mux_inst_897 (
  .O(mux_o_897),
  .I0(mux_o_893),
  .I1(mux_o_894),
  .S0(dff_q_5)
);
MUX2 mux_inst_898 (
  .O(mux_o_898),
  .I0(mux_o_895),
  .I1(mux_o_896),
  .S0(dff_q_5)
);
MUX2 mux_inst_899 (
  .O(doutb[27]),
  .I0(mux_o_897),
  .I1(mux_o_898),
  .S0(dff_q_4)
);
MUX2 mux_inst_900 (
  .O(mux_o_900),
  .I0(dpb_inst_16_doutb[28]),
  .I1(dpb_inst_17_doutb[28]),
  .S0(dff_q_7)
);
MUX2 mux_inst_901 (
  .O(mux_o_901),
  .I0(dpb_inst_18_doutb[28]),
  .I1(dpb_inst_19_doutb[28]),
  .S0(dff_q_7)
);
MUX2 mux_inst_902 (
  .O(mux_o_902),
  .I0(dpb_inst_20_doutb[28]),
  .I1(dpb_inst_21_doutb[28]),
  .S0(dff_q_7)
);
MUX2 mux_inst_903 (
  .O(mux_o_903),
  .I0(dpb_inst_22_doutb[28]),
  .I1(dpb_inst_23_doutb[28]),
  .S0(dff_q_7)
);
MUX2 mux_inst_904 (
  .O(mux_o_904),
  .I0(dpb_inst_24_doutb[28]),
  .I1(dpb_inst_25_doutb[28]),
  .S0(dff_q_7)
);
MUX2 mux_inst_905 (
  .O(mux_o_905),
  .I0(dpb_inst_26_doutb[28]),
  .I1(dpb_inst_27_doutb[28]),
  .S0(dff_q_7)
);
MUX2 mux_inst_906 (
  .O(mux_o_906),
  .I0(dpb_inst_28_doutb[28]),
  .I1(dpb_inst_29_doutb[28]),
  .S0(dff_q_7)
);
MUX2 mux_inst_907 (
  .O(mux_o_907),
  .I0(dpb_inst_30_doutb[28]),
  .I1(dpb_inst_31_doutb[28]),
  .S0(dff_q_7)
);
MUX2 mux_inst_908 (
  .O(mux_o_908),
  .I0(mux_o_900),
  .I1(mux_o_901),
  .S0(dff_q_6)
);
MUX2 mux_inst_909 (
  .O(mux_o_909),
  .I0(mux_o_902),
  .I1(mux_o_903),
  .S0(dff_q_6)
);
MUX2 mux_inst_910 (
  .O(mux_o_910),
  .I0(mux_o_904),
  .I1(mux_o_905),
  .S0(dff_q_6)
);
MUX2 mux_inst_911 (
  .O(mux_o_911),
  .I0(mux_o_906),
  .I1(mux_o_907),
  .S0(dff_q_6)
);
MUX2 mux_inst_912 (
  .O(mux_o_912),
  .I0(mux_o_908),
  .I1(mux_o_909),
  .S0(dff_q_5)
);
MUX2 mux_inst_913 (
  .O(mux_o_913),
  .I0(mux_o_910),
  .I1(mux_o_911),
  .S0(dff_q_5)
);
MUX2 mux_inst_914 (
  .O(doutb[28]),
  .I0(mux_o_912),
  .I1(mux_o_913),
  .S0(dff_q_4)
);
MUX2 mux_inst_915 (
  .O(mux_o_915),
  .I0(dpb_inst_16_doutb[29]),
  .I1(dpb_inst_17_doutb[29]),
  .S0(dff_q_7)
);
MUX2 mux_inst_916 (
  .O(mux_o_916),
  .I0(dpb_inst_18_doutb[29]),
  .I1(dpb_inst_19_doutb[29]),
  .S0(dff_q_7)
);
MUX2 mux_inst_917 (
  .O(mux_o_917),
  .I0(dpb_inst_20_doutb[29]),
  .I1(dpb_inst_21_doutb[29]),
  .S0(dff_q_7)
);
MUX2 mux_inst_918 (
  .O(mux_o_918),
  .I0(dpb_inst_22_doutb[29]),
  .I1(dpb_inst_23_doutb[29]),
  .S0(dff_q_7)
);
MUX2 mux_inst_919 (
  .O(mux_o_919),
  .I0(dpb_inst_24_doutb[29]),
  .I1(dpb_inst_25_doutb[29]),
  .S0(dff_q_7)
);
MUX2 mux_inst_920 (
  .O(mux_o_920),
  .I0(dpb_inst_26_doutb[29]),
  .I1(dpb_inst_27_doutb[29]),
  .S0(dff_q_7)
);
MUX2 mux_inst_921 (
  .O(mux_o_921),
  .I0(dpb_inst_28_doutb[29]),
  .I1(dpb_inst_29_doutb[29]),
  .S0(dff_q_7)
);
MUX2 mux_inst_922 (
  .O(mux_o_922),
  .I0(dpb_inst_30_doutb[29]),
  .I1(dpb_inst_31_doutb[29]),
  .S0(dff_q_7)
);
MUX2 mux_inst_923 (
  .O(mux_o_923),
  .I0(mux_o_915),
  .I1(mux_o_916),
  .S0(dff_q_6)
);
MUX2 mux_inst_924 (
  .O(mux_o_924),
  .I0(mux_o_917),
  .I1(mux_o_918),
  .S0(dff_q_6)
);
MUX2 mux_inst_925 (
  .O(mux_o_925),
  .I0(mux_o_919),
  .I1(mux_o_920),
  .S0(dff_q_6)
);
MUX2 mux_inst_926 (
  .O(mux_o_926),
  .I0(mux_o_921),
  .I1(mux_o_922),
  .S0(dff_q_6)
);
MUX2 mux_inst_927 (
  .O(mux_o_927),
  .I0(mux_o_923),
  .I1(mux_o_924),
  .S0(dff_q_5)
);
MUX2 mux_inst_928 (
  .O(mux_o_928),
  .I0(mux_o_925),
  .I1(mux_o_926),
  .S0(dff_q_5)
);
MUX2 mux_inst_929 (
  .O(doutb[29]),
  .I0(mux_o_927),
  .I1(mux_o_928),
  .S0(dff_q_4)
);
MUX2 mux_inst_930 (
  .O(mux_o_930),
  .I0(dpb_inst_16_doutb[30]),
  .I1(dpb_inst_17_doutb[30]),
  .S0(dff_q_7)
);
MUX2 mux_inst_931 (
  .O(mux_o_931),
  .I0(dpb_inst_18_doutb[30]),
  .I1(dpb_inst_19_doutb[30]),
  .S0(dff_q_7)
);
MUX2 mux_inst_932 (
  .O(mux_o_932),
  .I0(dpb_inst_20_doutb[30]),
  .I1(dpb_inst_21_doutb[30]),
  .S0(dff_q_7)
);
MUX2 mux_inst_933 (
  .O(mux_o_933),
  .I0(dpb_inst_22_doutb[30]),
  .I1(dpb_inst_23_doutb[30]),
  .S0(dff_q_7)
);
MUX2 mux_inst_934 (
  .O(mux_o_934),
  .I0(dpb_inst_24_doutb[30]),
  .I1(dpb_inst_25_doutb[30]),
  .S0(dff_q_7)
);
MUX2 mux_inst_935 (
  .O(mux_o_935),
  .I0(dpb_inst_26_doutb[30]),
  .I1(dpb_inst_27_doutb[30]),
  .S0(dff_q_7)
);
MUX2 mux_inst_936 (
  .O(mux_o_936),
  .I0(dpb_inst_28_doutb[30]),
  .I1(dpb_inst_29_doutb[30]),
  .S0(dff_q_7)
);
MUX2 mux_inst_937 (
  .O(mux_o_937),
  .I0(dpb_inst_30_doutb[30]),
  .I1(dpb_inst_31_doutb[30]),
  .S0(dff_q_7)
);
MUX2 mux_inst_938 (
  .O(mux_o_938),
  .I0(mux_o_930),
  .I1(mux_o_931),
  .S0(dff_q_6)
);
MUX2 mux_inst_939 (
  .O(mux_o_939),
  .I0(mux_o_932),
  .I1(mux_o_933),
  .S0(dff_q_6)
);
MUX2 mux_inst_940 (
  .O(mux_o_940),
  .I0(mux_o_934),
  .I1(mux_o_935),
  .S0(dff_q_6)
);
MUX2 mux_inst_941 (
  .O(mux_o_941),
  .I0(mux_o_936),
  .I1(mux_o_937),
  .S0(dff_q_6)
);
MUX2 mux_inst_942 (
  .O(mux_o_942),
  .I0(mux_o_938),
  .I1(mux_o_939),
  .S0(dff_q_5)
);
MUX2 mux_inst_943 (
  .O(mux_o_943),
  .I0(mux_o_940),
  .I1(mux_o_941),
  .S0(dff_q_5)
);
MUX2 mux_inst_944 (
  .O(doutb[30]),
  .I0(mux_o_942),
  .I1(mux_o_943),
  .S0(dff_q_4)
);
MUX2 mux_inst_945 (
  .O(mux_o_945),
  .I0(dpb_inst_16_doutb[31]),
  .I1(dpb_inst_17_doutb[31]),
  .S0(dff_q_7)
);
MUX2 mux_inst_946 (
  .O(mux_o_946),
  .I0(dpb_inst_18_doutb[31]),
  .I1(dpb_inst_19_doutb[31]),
  .S0(dff_q_7)
);
MUX2 mux_inst_947 (
  .O(mux_o_947),
  .I0(dpb_inst_20_doutb[31]),
  .I1(dpb_inst_21_doutb[31]),
  .S0(dff_q_7)
);
MUX2 mux_inst_948 (
  .O(mux_o_948),
  .I0(dpb_inst_22_doutb[31]),
  .I1(dpb_inst_23_doutb[31]),
  .S0(dff_q_7)
);
MUX2 mux_inst_949 (
  .O(mux_o_949),
  .I0(dpb_inst_24_doutb[31]),
  .I1(dpb_inst_25_doutb[31]),
  .S0(dff_q_7)
);
MUX2 mux_inst_950 (
  .O(mux_o_950),
  .I0(dpb_inst_26_doutb[31]),
  .I1(dpb_inst_27_doutb[31]),
  .S0(dff_q_7)
);
MUX2 mux_inst_951 (
  .O(mux_o_951),
  .I0(dpb_inst_28_doutb[31]),
  .I1(dpb_inst_29_doutb[31]),
  .S0(dff_q_7)
);
MUX2 mux_inst_952 (
  .O(mux_o_952),
  .I0(dpb_inst_30_doutb[31]),
  .I1(dpb_inst_31_doutb[31]),
  .S0(dff_q_7)
);
MUX2 mux_inst_953 (
  .O(mux_o_953),
  .I0(mux_o_945),
  .I1(mux_o_946),
  .S0(dff_q_6)
);
MUX2 mux_inst_954 (
  .O(mux_o_954),
  .I0(mux_o_947),
  .I1(mux_o_948),
  .S0(dff_q_6)
);
MUX2 mux_inst_955 (
  .O(mux_o_955),
  .I0(mux_o_949),
  .I1(mux_o_950),
  .S0(dff_q_6)
);
MUX2 mux_inst_956 (
  .O(mux_o_956),
  .I0(mux_o_951),
  .I1(mux_o_952),
  .S0(dff_q_6)
);
MUX2 mux_inst_957 (
  .O(mux_o_957),
  .I0(mux_o_953),
  .I1(mux_o_954),
  .S0(dff_q_5)
);
MUX2 mux_inst_958 (
  .O(mux_o_958),
  .I0(mux_o_955),
  .I1(mux_o_956),
  .S0(dff_q_5)
);
MUX2 mux_inst_959 (
  .O(doutb[31]),
  .I0(mux_o_957),
  .I1(mux_o_958),
  .S0(dff_q_4)
);
endmodule //Gowin_DPB
