TORVS/torvs9p1.sv