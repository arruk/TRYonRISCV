TORVS/torvs5C.sv