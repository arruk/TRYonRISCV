//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.10.03 Education
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Device Version: C
//Created Time: Fri Jan 10 18:43:48 2025

module Gowin_DPB (douta, doutb, clka, ocea, cea, reseta, wrea, clkb, oceb, ceb, resetb, wreb, ada, dina, adb, dinb, byte_ena, byte_enb);

output [31:0] douta;
output [31:0] doutb;
input clka;
input ocea;
input cea;
input reseta;
input wrea;
input clkb;
input oceb;
input ceb;
input resetb;
input wreb;
input [13:0] ada;
input [31:0] dina;
input [13:0] adb;
input [31:0] dinb;
input [3:0] byte_ena;
input [3:0] byte_enb;

wire [8:0] dpx9b_inst_0_douta_w;
wire [8:0] dpx9b_inst_0_douta;
wire [8:0] dpx9b_inst_0_doutb_w;
wire [8:0] dpx9b_inst_0_doutb;
wire [8:0] dpx9b_inst_1_douta_w;
wire [8:0] dpx9b_inst_1_douta;
wire [8:0] dpx9b_inst_1_doutb_w;
wire [8:0] dpx9b_inst_1_doutb;
wire [8:0] dpx9b_inst_2_douta_w;
wire [8:0] dpx9b_inst_2_douta;
wire [8:0] dpx9b_inst_2_doutb_w;
wire [8:0] dpx9b_inst_2_doutb;
wire [8:0] dpx9b_inst_3_douta_w;
wire [8:0] dpx9b_inst_3_douta;
wire [8:0] dpx9b_inst_3_doutb_w;
wire [8:0] dpx9b_inst_3_doutb;
wire [8:0] dpx9b_inst_4_douta_w;
wire [8:0] dpx9b_inst_4_douta;
wire [8:0] dpx9b_inst_4_doutb_w;
wire [8:0] dpx9b_inst_4_doutb;
wire [8:0] dpx9b_inst_5_douta_w;
wire [8:0] dpx9b_inst_5_douta;
wire [8:0] dpx9b_inst_5_doutb_w;
wire [8:0] dpx9b_inst_5_doutb;
wire [8:0] dpx9b_inst_6_douta_w;
wire [8:0] dpx9b_inst_6_douta;
wire [8:0] dpx9b_inst_6_doutb_w;
wire [8:0] dpx9b_inst_6_doutb;
wire [8:0] dpx9b_inst_7_douta_w;
wire [8:0] dpx9b_inst_7_douta;
wire [8:0] dpx9b_inst_7_doutb_w;
wire [8:0] dpx9b_inst_7_doutb;
wire [8:0] dpx9b_inst_8_douta_w;
wire [17:9] dpx9b_inst_8_douta;
wire [8:0] dpx9b_inst_8_doutb_w;
wire [17:9] dpx9b_inst_8_doutb;
wire [8:0] dpx9b_inst_9_douta_w;
wire [17:9] dpx9b_inst_9_douta;
wire [8:0] dpx9b_inst_9_doutb_w;
wire [17:9] dpx9b_inst_9_doutb;
wire [8:0] dpx9b_inst_10_douta_w;
wire [17:9] dpx9b_inst_10_douta;
wire [8:0] dpx9b_inst_10_doutb_w;
wire [17:9] dpx9b_inst_10_doutb;
wire [8:0] dpx9b_inst_11_douta_w;
wire [17:9] dpx9b_inst_11_douta;
wire [8:0] dpx9b_inst_11_doutb_w;
wire [17:9] dpx9b_inst_11_doutb;
wire [8:0] dpx9b_inst_12_douta_w;
wire [17:9] dpx9b_inst_12_douta;
wire [8:0] dpx9b_inst_12_doutb_w;
wire [17:9] dpx9b_inst_12_doutb;
wire [8:0] dpx9b_inst_13_douta_w;
wire [17:9] dpx9b_inst_13_douta;
wire [8:0] dpx9b_inst_13_doutb_w;
wire [17:9] dpx9b_inst_13_doutb;
wire [8:0] dpx9b_inst_14_douta_w;
wire [17:9] dpx9b_inst_14_douta;
wire [8:0] dpx9b_inst_14_doutb_w;
wire [17:9] dpx9b_inst_14_doutb;
wire [8:0] dpx9b_inst_15_douta_w;
wire [17:9] dpx9b_inst_15_douta;
wire [8:0] dpx9b_inst_15_doutb_w;
wire [17:9] dpx9b_inst_15_doutb;
wire [8:0] dpx9b_inst_16_douta_w;
wire [26:18] dpx9b_inst_16_douta;
wire [8:0] dpx9b_inst_16_doutb_w;
wire [26:18] dpx9b_inst_16_doutb;
wire [8:0] dpx9b_inst_17_douta_w;
wire [26:18] dpx9b_inst_17_douta;
wire [8:0] dpx9b_inst_17_doutb_w;
wire [26:18] dpx9b_inst_17_doutb;
wire [8:0] dpx9b_inst_18_douta_w;
wire [26:18] dpx9b_inst_18_douta;
wire [8:0] dpx9b_inst_18_doutb_w;
wire [26:18] dpx9b_inst_18_doutb;
wire [8:0] dpx9b_inst_19_douta_w;
wire [26:18] dpx9b_inst_19_douta;
wire [8:0] dpx9b_inst_19_doutb_w;
wire [26:18] dpx9b_inst_19_doutb;
wire [8:0] dpx9b_inst_20_douta_w;
wire [26:18] dpx9b_inst_20_douta;
wire [8:0] dpx9b_inst_20_doutb_w;
wire [26:18] dpx9b_inst_20_doutb;
wire [8:0] dpx9b_inst_21_douta_w;
wire [26:18] dpx9b_inst_21_douta;
wire [8:0] dpx9b_inst_21_doutb_w;
wire [26:18] dpx9b_inst_21_doutb;
wire [8:0] dpx9b_inst_22_douta_w;
wire [26:18] dpx9b_inst_22_douta;
wire [8:0] dpx9b_inst_22_doutb_w;
wire [26:18] dpx9b_inst_22_doutb;
wire [8:0] dpx9b_inst_23_douta_w;
wire [26:18] dpx9b_inst_23_douta;
wire [8:0] dpx9b_inst_23_doutb_w;
wire [26:18] dpx9b_inst_23_doutb;
wire [14:0] dpb_inst_24_douta_w;
wire [14:0] dpb_inst_24_doutb_w;
wire [14:0] dpb_inst_25_douta_w;
wire [14:0] dpb_inst_25_doutb_w;
wire [14:0] dpb_inst_26_douta_w;
wire [14:0] dpb_inst_26_doutb_w;
wire [14:0] dpb_inst_27_douta_w;
wire [14:0] dpb_inst_27_doutb_w;
wire [14:0] dpb_inst_28_douta_w;
wire [14:0] dpb_inst_28_doutb_w;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire dff_q_4;
wire dff_q_5;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;
wire mux_o_7;
wire mux_o_8;
wire mux_o_9;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_14;
wire mux_o_15;
wire mux_o_16;
wire mux_o_17;
wire mux_o_18;
wire mux_o_19;
wire mux_o_21;
wire mux_o_22;
wire mux_o_23;
wire mux_o_24;
wire mux_o_25;
wire mux_o_26;
wire mux_o_28;
wire mux_o_29;
wire mux_o_30;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_35;
wire mux_o_36;
wire mux_o_37;
wire mux_o_38;
wire mux_o_39;
wire mux_o_40;
wire mux_o_42;
wire mux_o_43;
wire mux_o_44;
wire mux_o_45;
wire mux_o_46;
wire mux_o_47;
wire mux_o_49;
wire mux_o_50;
wire mux_o_51;
wire mux_o_52;
wire mux_o_53;
wire mux_o_54;
wire mux_o_56;
wire mux_o_57;
wire mux_o_58;
wire mux_o_59;
wire mux_o_60;
wire mux_o_61;
wire mux_o_63;
wire mux_o_64;
wire mux_o_65;
wire mux_o_66;
wire mux_o_67;
wire mux_o_68;
wire mux_o_70;
wire mux_o_71;
wire mux_o_72;
wire mux_o_73;
wire mux_o_74;
wire mux_o_75;
wire mux_o_77;
wire mux_o_78;
wire mux_o_79;
wire mux_o_80;
wire mux_o_81;
wire mux_o_82;
wire mux_o_84;
wire mux_o_85;
wire mux_o_86;
wire mux_o_87;
wire mux_o_88;
wire mux_o_89;
wire mux_o_91;
wire mux_o_92;
wire mux_o_93;
wire mux_o_94;
wire mux_o_95;
wire mux_o_96;
wire mux_o_98;
wire mux_o_99;
wire mux_o_100;
wire mux_o_101;
wire mux_o_102;
wire mux_o_103;
wire mux_o_105;
wire mux_o_106;
wire mux_o_107;
wire mux_o_108;
wire mux_o_109;
wire mux_o_110;
wire mux_o_112;
wire mux_o_113;
wire mux_o_114;
wire mux_o_115;
wire mux_o_116;
wire mux_o_117;
wire mux_o_119;
wire mux_o_120;
wire mux_o_121;
wire mux_o_122;
wire mux_o_123;
wire mux_o_124;
wire mux_o_126;
wire mux_o_127;
wire mux_o_128;
wire mux_o_129;
wire mux_o_130;
wire mux_o_131;
wire mux_o_133;
wire mux_o_134;
wire mux_o_135;
wire mux_o_136;
wire mux_o_137;
wire mux_o_138;
wire mux_o_140;
wire mux_o_141;
wire mux_o_142;
wire mux_o_143;
wire mux_o_144;
wire mux_o_145;
wire mux_o_147;
wire mux_o_148;
wire mux_o_149;
wire mux_o_150;
wire mux_o_151;
wire mux_o_152;
wire mux_o_154;
wire mux_o_155;
wire mux_o_156;
wire mux_o_157;
wire mux_o_158;
wire mux_o_159;
wire mux_o_161;
wire mux_o_162;
wire mux_o_163;
wire mux_o_164;
wire mux_o_165;
wire mux_o_166;
wire mux_o_168;
wire mux_o_169;
wire mux_o_170;
wire mux_o_171;
wire mux_o_172;
wire mux_o_173;
wire mux_o_175;
wire mux_o_176;
wire mux_o_177;
wire mux_o_178;
wire mux_o_179;
wire mux_o_180;
wire mux_o_182;
wire mux_o_183;
wire mux_o_184;
wire mux_o_185;
wire mux_o_186;
wire mux_o_187;
wire mux_o_189;
wire mux_o_190;
wire mux_o_191;
wire mux_o_192;
wire mux_o_193;
wire mux_o_194;
wire mux_o_196;
wire mux_o_197;
wire mux_o_198;
wire mux_o_199;
wire mux_o_200;
wire mux_o_201;
wire mux_o_203;
wire mux_o_204;
wire mux_o_205;
wire mux_o_206;
wire mux_o_207;
wire mux_o_208;
wire mux_o_210;
wire mux_o_211;
wire mux_o_212;
wire mux_o_213;
wire mux_o_214;
wire mux_o_215;
wire mux_o_217;
wire mux_o_218;
wire mux_o_219;
wire mux_o_220;
wire mux_o_221;
wire mux_o_222;
wire mux_o_224;
wire mux_o_225;
wire mux_o_226;
wire mux_o_227;
wire mux_o_228;
wire mux_o_229;
wire mux_o_231;
wire mux_o_232;
wire mux_o_233;
wire mux_o_234;
wire mux_o_235;
wire mux_o_236;
wire mux_o_238;
wire mux_o_239;
wire mux_o_240;
wire mux_o_241;
wire mux_o_242;
wire mux_o_243;
wire mux_o_245;
wire mux_o_246;
wire mux_o_247;
wire mux_o_248;
wire mux_o_249;
wire mux_o_250;
wire mux_o_252;
wire mux_o_253;
wire mux_o_254;
wire mux_o_255;
wire mux_o_256;
wire mux_o_257;
wire mux_o_259;
wire mux_o_260;
wire mux_o_261;
wire mux_o_262;
wire mux_o_263;
wire mux_o_264;
wire mux_o_266;
wire mux_o_267;
wire mux_o_268;
wire mux_o_269;
wire mux_o_270;
wire mux_o_271;
wire mux_o_273;
wire mux_o_274;
wire mux_o_275;
wire mux_o_276;
wire mux_o_277;
wire mux_o_278;
wire mux_o_280;
wire mux_o_281;
wire mux_o_282;
wire mux_o_283;
wire mux_o_284;
wire mux_o_285;
wire mux_o_287;
wire mux_o_288;
wire mux_o_289;
wire mux_o_290;
wire mux_o_291;
wire mux_o_292;
wire mux_o_294;
wire mux_o_295;
wire mux_o_296;
wire mux_o_297;
wire mux_o_298;
wire mux_o_299;
wire mux_o_301;
wire mux_o_302;
wire mux_o_303;
wire mux_o_304;
wire mux_o_305;
wire mux_o_306;
wire mux_o_308;
wire mux_o_309;
wire mux_o_310;
wire mux_o_311;
wire mux_o_312;
wire mux_o_313;
wire mux_o_315;
wire mux_o_316;
wire mux_o_317;
wire mux_o_318;
wire mux_o_319;
wire mux_o_320;
wire mux_o_322;
wire mux_o_323;
wire mux_o_324;
wire mux_o_325;
wire mux_o_326;
wire mux_o_327;
wire mux_o_329;
wire mux_o_330;
wire mux_o_331;
wire mux_o_332;
wire mux_o_333;
wire mux_o_334;
wire mux_o_336;
wire mux_o_337;
wire mux_o_338;
wire mux_o_339;
wire mux_o_340;
wire mux_o_341;
wire mux_o_343;
wire mux_o_344;
wire mux_o_345;
wire mux_o_346;
wire mux_o_347;
wire mux_o_348;
wire mux_o_350;
wire mux_o_351;
wire mux_o_352;
wire mux_o_353;
wire mux_o_354;
wire mux_o_355;
wire mux_o_357;
wire mux_o_358;
wire mux_o_359;
wire mux_o_360;
wire mux_o_361;
wire mux_o_362;
wire mux_o_364;
wire mux_o_365;
wire mux_o_366;
wire mux_o_367;
wire mux_o_368;
wire mux_o_369;
wire mux_o_371;
wire mux_o_372;
wire mux_o_373;
wire mux_o_374;
wire mux_o_375;
wire mux_o_376;
wire cea_w;
wire ceb_w;
wire gw_gnd;

assign cea_w = ~wrea & cea;
assign ceb_w = ~wreb & ceb;
assign gw_gnd = 1'b0;

DPX9B dpx9b_inst_0 (
    .DOA({dpx9b_inst_0_douta_w[8:0],dpx9b_inst_0_douta[8:0]}),
    .DOB({dpx9b_inst_0_doutb_w[8:0],dpx9b_inst_0_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_0.READ_MODE0 = 1'b0;
defparam dpx9b_inst_0.READ_MODE1 = 1'b0;
defparam dpx9b_inst_0.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_0.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_0.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_0.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_0.BLK_SEL_0 = 3'b000;
defparam dpx9b_inst_0.BLK_SEL_1 = 3'b000;
defparam dpx9b_inst_0.RESET_MODE = "SYNC";
defparam dpx9b_inst_0.INIT_RAM_00 = 288'h10082E62030DB8CA7322538A74F26D3C8A53220287B65B18F8143DB91A47C3D218F84A25;
defparam dpx9b_inst_0.INIT_RAM_01 = 288'h32DB8E869B9940CA6930996CF20B4480D363B9142E972905D2CA68901A6C7722850ECF6E;
defparam dpx9b_inst_0.INIT_RAM_02 = 288'h3A914C873B75087C64B6DBA843E001BEE468B91CC402C309B8EA451D5B4CB68339A2DC66;
defparam dpx9b_inst_0.INIT_RAM_03 = 288'hAFD080120329B0E620100024020100E88E4900186DC6537194E661BB1D2416C3651AC86E;
defparam dpx9b_inst_0.INIT_RAM_04 = 288'h90080BA6F98904012010080C55F218024065361CC40200048040203157C8600900804062;
defparam dpx9b_inst_0.INIT_RAM_05 = 288'h39880400090080406DB90805A4728000567527D884065361CC402000480755D37CC88200;
defparam dpx9b_inst_0.INIT_RAM_06 = 288'hB9080012010080DB74100024020105BEEA20004804020105CC406E328B6E86538080CA6C;
defparam dpx9b_inst_0.INIT_RAM_07 = 288'h16DD0CA7010194D87310082C55F2FD389320A9D06A54EAC880CA6C39880400090080406D;
defparam dpx9b_inst_0.INIT_RAM_08 = 288'h10080745F2280240201018E664900480402031CC8920090080406398926ED2032C80DC65;
defparam dpx9b_inst_0.INIT_RAM_09 = 288'h3988040009008040639914C932098D06A54EAC880CA6C3988040009008040639894C0120;
defparam dpx9b_inst_0.INIT_RAM_0A = 288'h325904A6FBADB8CB65A19BA402C31990CA5FAA896DD6632D38932099506A54EAC880CA6C;
defparam dpx9b_inst_0.INIT_RAM_0B = 288'hA714C4E4DA7914A644A714E4E4DA7914A64405094C87AB954E88643D5CAC96532D94E644;
defparam dpx9b_inst_0.INIT_RAM_0C = 288'h83C1E0E06030180C06030180D0582C160A040240E000021CE26930A714C4E4DA7914A644;
defparam dpx9b_inst_0.INIT_RAM_0D = 288'h04020100804020100804020100804020100804020110783C1E0F0783C1E0F0783C1E0F07;
defparam dpx9b_inst_0.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000008040201008040201008040201008;
defparam dpx9b_inst_0.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_0.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_1 (
    .DOA({dpx9b_inst_1_douta_w[8:0],dpx9b_inst_1_douta[8:0]}),
    .DOB({dpx9b_inst_1_doutb_w[8:0],dpx9b_inst_1_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_1.READ_MODE0 = 1'b0;
defparam dpx9b_inst_1.READ_MODE1 = 1'b0;
defparam dpx9b_inst_1.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_1.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_1.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_1.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_1.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_1.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_1.RESET_MODE = "SYNC";
defparam dpx9b_inst_1.INIT_RAM_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_1E = 288'hF6060A11B008040010000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_1F = 288'h8200411740052360182846C020100040164422110884422111710C854200B01821D0002C;
defparam dpx9b_inst_1.INIT_RAM_20 = 288'h2211088708541C0A02845B001D448060911B008040010059108844221108844B64321306;
defparam dpx9b_inst_1.INIT_RAM_21 = 288'h00000000B225128944A2512150C8541C0908819C000F002060991B008040010059108844;
defparam dpx9b_inst_1.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_1.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_2 (
    .DOA({dpx9b_inst_2_douta_w[8:0],dpx9b_inst_2_douta[8:0]}),
    .DOB({dpx9b_inst_2_doutb_w[8:0],dpx9b_inst_2_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_2.READ_MODE0 = 1'b0;
defparam dpx9b_inst_2.READ_MODE1 = 1'b0;
defparam dpx9b_inst_2.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_2.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_2.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_2.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_2.BLK_SEL_0 = 3'b010;
defparam dpx9b_inst_2.BLK_SEL_1 = 3'b010;
defparam dpx9b_inst_2.RESET_MODE = "SYNC";
defparam dpx9b_inst_2.INIT_RAM_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_2.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_3 (
    .DOA({dpx9b_inst_3_douta_w[8:0],dpx9b_inst_3_douta[8:0]}),
    .DOB({dpx9b_inst_3_doutb_w[8:0],dpx9b_inst_3_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_3.READ_MODE0 = 1'b0;
defparam dpx9b_inst_3.READ_MODE1 = 1'b0;
defparam dpx9b_inst_3.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_3.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_3.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_3.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_3.BLK_SEL_0 = 3'b011;
defparam dpx9b_inst_3.BLK_SEL_1 = 3'b011;
defparam dpx9b_inst_3.RESET_MODE = "SYNC";
defparam dpx9b_inst_3.INIT_RAM_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_3.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_4 (
    .DOA({dpx9b_inst_4_douta_w[8:0],dpx9b_inst_4_douta[8:0]}),
    .DOB({dpx9b_inst_4_doutb_w[8:0],dpx9b_inst_4_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_4.READ_MODE0 = 1'b0;
defparam dpx9b_inst_4.READ_MODE1 = 1'b0;
defparam dpx9b_inst_4.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_4.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_4.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_4.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_4.BLK_SEL_0 = 3'b100;
defparam dpx9b_inst_4.BLK_SEL_1 = 3'b100;
defparam dpx9b_inst_4.RESET_MODE = "SYNC";
defparam dpx9b_inst_4.INIT_RAM_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_4.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_5 (
    .DOA({dpx9b_inst_5_douta_w[8:0],dpx9b_inst_5_douta[8:0]}),
    .DOB({dpx9b_inst_5_doutb_w[8:0],dpx9b_inst_5_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_5.READ_MODE0 = 1'b0;
defparam dpx9b_inst_5.READ_MODE1 = 1'b0;
defparam dpx9b_inst_5.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_5.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_5.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_5.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_5.BLK_SEL_0 = 3'b101;
defparam dpx9b_inst_5.BLK_SEL_1 = 3'b101;
defparam dpx9b_inst_5.RESET_MODE = "SYNC";
defparam dpx9b_inst_5.INIT_RAM_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_5.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_6 (
    .DOA({dpx9b_inst_6_douta_w[8:0],dpx9b_inst_6_douta[8:0]}),
    .DOB({dpx9b_inst_6_doutb_w[8:0],dpx9b_inst_6_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_6.READ_MODE0 = 1'b0;
defparam dpx9b_inst_6.READ_MODE1 = 1'b0;
defparam dpx9b_inst_6.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_6.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_6.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_6.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_6.BLK_SEL_0 = 3'b110;
defparam dpx9b_inst_6.BLK_SEL_1 = 3'b110;
defparam dpx9b_inst_6.RESET_MODE = "SYNC";
defparam dpx9b_inst_6.INIT_RAM_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_6.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_7 (
    .DOA({dpx9b_inst_7_douta_w[8:0],dpx9b_inst_7_douta[8:0]}),
    .DOB({dpx9b_inst_7_doutb_w[8:0],dpx9b_inst_7_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_7.READ_MODE0 = 1'b0;
defparam dpx9b_inst_7.READ_MODE1 = 1'b0;
defparam dpx9b_inst_7.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_7.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_7.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_7.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_7.BLK_SEL_0 = 3'b111;
defparam dpx9b_inst_7.BLK_SEL_1 = 3'b111;
defparam dpx9b_inst_7.RESET_MODE = "SYNC";
defparam dpx9b_inst_7.INIT_RAM_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_7.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_8 (
    .DOA({dpx9b_inst_8_douta_w[8:0],dpx9b_inst_8_douta[17:9]}),
    .DOB({dpx9b_inst_8_doutb_w[8:0],dpx9b_inst_8_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_8.READ_MODE0 = 1'b0;
defparam dpx9b_inst_8.READ_MODE1 = 1'b0;
defparam dpx9b_inst_8.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_8.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_8.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_8.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_8.BLK_SEL_0 = 3'b000;
defparam dpx9b_inst_8.BLK_SEL_1 = 3'b000;
defparam dpx9b_inst_8.RESET_MODE = "SYNC";
defparam dpx9b_inst_8.INIT_RAM_00 = 288'h0A46768ABDC8C621BA9A08E54A60B48C21AA920012039DE47C0090196DE3E005447C6532;
defparam dpx9b_inst_8.INIT_RAM_01 = 288'h1CAE968BB192D800B11D6E769135BAED6CB7586E46534184C967905DAD96EB0DC85264B3;
defparam dpx9b_inst_8.INIT_RAM_02 = 288'h5D2F00AB757ECA3E05590BF651F002DF78105B84172901CE4174BC084C36E321A6E47310;
defparam dpx9b_inst_8.INIT_RAM_03 = 288'h11EDC00120E8CB6810080002410080436C37006E46310080C92031982D26EBA884D07290;
defparam dpx9b_inst_8.INIT_RAM_04 = 288'h090403BB1D7CE40192080403A23DA003241D196D020100064820100E88F680009040201D;
defparam dpx9b_inst_8.INIT_RAM_05 = 288'hDA0402000090402138D78403FB69D00121B7D9CC94E1D196D020100004821ADD8EBE7200;
defparam dpx9b_inst_8.INIT_RAM_06 = 288'hD7E4000120804271AF480002410080DB6C90000482010084C420BA1BACB68375B2503A32;
defparam dpx9b_inst_8.INIT_RAM_07 = 288'h596D06EB64A07465B4080422C23140CB4E295389B4E22148883A32DA0402000C90402138;
defparam dpx9b_inst_8.INIT_RAM_08 = 288'h0804021A65B8002410080745E370004820100E8BC6E0009040201D178DC6530482E57437;
defparam dpx9b_inst_8.INIT_RAM_09 = 288'hDA0402000C9040201D17CEB4E29C989B4E22148883A32DA0402000C9040201D17CE80012;
defparam dpx9b_inst_8.INIT_RAM_0A = 288'h0284A6537188E773B9DE01668905B6403AAA5CCCA732FDCAEB4E298989B4E22148883A32;
defparam dpx9b_inst_8.INIT_RAM_0B = 288'h11CA84E1691843552411CA85216918435524002C92E1D578BD4C050EABC5FB1DCEE77534;
defparam dpx9b_inst_8.INIT_RAM_0C = 288'hC1E0F070381C0E070381C0E068241209040201606000051272351811CA85216918435524;
defparam dpx9b_inst_8.INIT_RAM_0D = 288'h020100804020100804020100804020100804020100983C1E0F0783C1E0F0783C1E0F0783;
defparam dpx9b_inst_8.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000004020100804020100804020100804;
defparam dpx9b_inst_8.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_8.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_9 (
    .DOA({dpx9b_inst_9_douta_w[8:0],dpx9b_inst_9_douta[17:9]}),
    .DOB({dpx9b_inst_9_doutb_w[8:0],dpx9b_inst_9_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_9.READ_MODE0 = 1'b0;
defparam dpx9b_inst_9.READ_MODE1 = 1'b0;
defparam dpx9b_inst_9.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_9.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_9.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_9.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_9.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_9.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_9.RESET_MODE = "SYNC";
defparam dpx9b_inst_9.INIT_RAM_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_1E = 288'hB880001065F4F40000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_1F = 288'h64D1299C49100AE800004197D3D000000007369B0D66A3499202CDE632E95C4E55124403;
defparam dpx9b_inst_9.INIT_RAM_20 = 288'h351A4C901E632E9449607124402BB80001065F4F400000001CDA6C359A8D2648033799CA;
defparam dpx9b_inst_9.INIT_RAM_21 = 288'h000000000039B0D66A34990C001E632E94C064D124402BD00001065F4F400000001CD86B;
defparam dpx9b_inst_9.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_9.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_10 (
    .DOA({dpx9b_inst_10_douta_w[8:0],dpx9b_inst_10_douta[17:9]}),
    .DOB({dpx9b_inst_10_doutb_w[8:0],dpx9b_inst_10_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_10.READ_MODE0 = 1'b0;
defparam dpx9b_inst_10.READ_MODE1 = 1'b0;
defparam dpx9b_inst_10.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_10.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_10.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_10.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_10.BLK_SEL_0 = 3'b010;
defparam dpx9b_inst_10.BLK_SEL_1 = 3'b010;
defparam dpx9b_inst_10.RESET_MODE = "SYNC";
defparam dpx9b_inst_10.INIT_RAM_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_10.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_11 (
    .DOA({dpx9b_inst_11_douta_w[8:0],dpx9b_inst_11_douta[17:9]}),
    .DOB({dpx9b_inst_11_doutb_w[8:0],dpx9b_inst_11_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_11.READ_MODE0 = 1'b0;
defparam dpx9b_inst_11.READ_MODE1 = 1'b0;
defparam dpx9b_inst_11.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_11.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_11.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_11.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_11.BLK_SEL_0 = 3'b011;
defparam dpx9b_inst_11.BLK_SEL_1 = 3'b011;
defparam dpx9b_inst_11.RESET_MODE = "SYNC";
defparam dpx9b_inst_11.INIT_RAM_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_11.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_12 (
    .DOA({dpx9b_inst_12_douta_w[8:0],dpx9b_inst_12_douta[17:9]}),
    .DOB({dpx9b_inst_12_doutb_w[8:0],dpx9b_inst_12_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_12.READ_MODE0 = 1'b0;
defparam dpx9b_inst_12.READ_MODE1 = 1'b0;
defparam dpx9b_inst_12.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_12.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_12.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_12.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_12.BLK_SEL_0 = 3'b100;
defparam dpx9b_inst_12.BLK_SEL_1 = 3'b100;
defparam dpx9b_inst_12.RESET_MODE = "SYNC";
defparam dpx9b_inst_12.INIT_RAM_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_12.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_13 (
    .DOA({dpx9b_inst_13_douta_w[8:0],dpx9b_inst_13_douta[17:9]}),
    .DOB({dpx9b_inst_13_doutb_w[8:0],dpx9b_inst_13_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_13.READ_MODE0 = 1'b0;
defparam dpx9b_inst_13.READ_MODE1 = 1'b0;
defparam dpx9b_inst_13.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_13.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_13.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_13.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_13.BLK_SEL_0 = 3'b101;
defparam dpx9b_inst_13.BLK_SEL_1 = 3'b101;
defparam dpx9b_inst_13.RESET_MODE = "SYNC";
defparam dpx9b_inst_13.INIT_RAM_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_13.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_14 (
    .DOA({dpx9b_inst_14_douta_w[8:0],dpx9b_inst_14_douta[17:9]}),
    .DOB({dpx9b_inst_14_doutb_w[8:0],dpx9b_inst_14_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_14.READ_MODE0 = 1'b0;
defparam dpx9b_inst_14.READ_MODE1 = 1'b0;
defparam dpx9b_inst_14.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_14.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_14.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_14.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_14.BLK_SEL_0 = 3'b110;
defparam dpx9b_inst_14.BLK_SEL_1 = 3'b110;
defparam dpx9b_inst_14.RESET_MODE = "SYNC";
defparam dpx9b_inst_14.INIT_RAM_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_14.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_15 (
    .DOA({dpx9b_inst_15_douta_w[8:0],dpx9b_inst_15_douta[17:9]}),
    .DOB({dpx9b_inst_15_doutb_w[8:0],dpx9b_inst_15_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_15.READ_MODE0 = 1'b0;
defparam dpx9b_inst_15.READ_MODE1 = 1'b0;
defparam dpx9b_inst_15.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_15.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_15.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_15.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_15.BLK_SEL_0 = 3'b111;
defparam dpx9b_inst_15.BLK_SEL_1 = 3'b111;
defparam dpx9b_inst_15.RESET_MODE = "SYNC";
defparam dpx9b_inst_15.INIT_RAM_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_15.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_16 (
    .DOA({dpx9b_inst_16_douta_w[8:0],dpx9b_inst_16_douta[26:18]}),
    .DOB({dpx9b_inst_16_doutb_w[8:0],dpx9b_inst_16_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_16.READ_MODE0 = 1'b0;
defparam dpx9b_inst_16.READ_MODE1 = 1'b0;
defparam dpx9b_inst_16.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_16.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_16.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_16.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_16.BLK_SEL_0 = 3'b000;
defparam dpx9b_inst_16.BLK_SEL_1 = 3'b000;
defparam dpx9b_inst_16.RESET_MODE = "SYNC";
defparam dpx9b_inst_16.INIT_RAM_00 = 288'h2992F36998D56AA19B2E000A8116415129932A00212088C03C01090EC701E000903C000B;
defparam dpx9b_inst_16.INIT_RAM_01 = 288'hE426C3219E4164011D4E826395C8EC6A321B0DF6C01588EF71B4898D464361BED8001C5D;
defparam dpx9b_inst_16.INIT_RAM_02 = 288'hED364014FCD1641E00A7974B20F002663811EE8773B096EC73B4D90037030888456E115C;
defparam dpx9b_inst_16.INIT_RAM_03 = 288'hEDC6C009904222B6080400132080402137DD0026AB5580E921BB5B2E06432D92E96C0199;
defparam dpx9b_inst_16.INIT_RAM_04 = 288'h4C820101688F7000980402011DB4B80130084456C10080026010080476CAE004C8201008;
defparam dpx9b_inst_16.INIT_RAM_05 = 288'hAD82010004C820100EE8450009BEE000181C4BF72BA084456C100800264114D0B447B800;
defparam dpx9b_inst_16.INIT_RAM_06 = 288'hE84500099040201DD0C9001320804271AF9100264100804270A20AAC867365DACD681088;
defparam dpx9b_inst_16.INIT_RAM_07 = 288'h0CE6CBB59AD021115B040201FDB4EC782295A982D2208EAA481088AD82010004E020100E;
defparam dpx9b_inst_16.INIT_RAM_08 = 288'h0402010DBAE801320804023A7DD0026410080474FBA004C8201008E9F7401D86C5621559;
defparam dpx9b_inst_16.INIT_RAM_09 = 288'hAD82010004E0201008E9F7022958A02D2208EAA481088AD82010004E0201008E9F700099;
defparam dpx9b_inst_16.INIT_RAM_0A = 288'h00566960E2EA74AE178C001B7096C962915A4C8081D54EBA6C22958982D2208EAA481088;
defparam dpx9b_inst_16.INIT_RAM_0B = 288'h0015022882A2532654001502A482A253265400426134809D502400A404EA99B6B85F365C;
defparam dpx9b_inst_16.INIT_RAM_0C = 288'hE0F078381C0E070381C0E070341A0D06830180B010000C8A439ACC0015022C82A2532654;
defparam dpx9b_inst_16.INIT_RAM_0D = 288'h0100804020100804020100804020100804020100805C1E0F0783C1E0F0783C1E0F0783C1;
defparam dpx9b_inst_16.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000002010080402010080402010080402;
defparam dpx9b_inst_16.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_16.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_17 (
    .DOA({dpx9b_inst_17_douta_w[8:0],dpx9b_inst_17_douta[26:18]}),
    .DOB({dpx9b_inst_17_doutb_w[8:0],dpx9b_inst_17_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_17.READ_MODE0 = 1'b0;
defparam dpx9b_inst_17.READ_MODE1 = 1'b0;
defparam dpx9b_inst_17.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_17.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_17.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_17.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_17.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_17.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_17.RESET_MODE = "SYNC";
defparam dpx9b_inst_17.INIT_RAM_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_1E = 288'hFF8000000200500000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_1F = 288'h80A00858001803FE0000000801400000010068947A3516894484C34100B02C020A000600;
defparam dpx9b_inst_17.INIT_RAM_20 = 288'hA8B44A2426100A82C1006000600FF800000020050000000401A251E8D45A2512130D05C1;
defparam dpx9b_inst_17.INIT_RAM_21 = 288'h00000000080244239188A4422484100A8280C09000600FF800000020050000000400A3D1;
defparam dpx9b_inst_17.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_17.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_18 (
    .DOA({dpx9b_inst_18_douta_w[8:0],dpx9b_inst_18_douta[26:18]}),
    .DOB({dpx9b_inst_18_doutb_w[8:0],dpx9b_inst_18_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_18.READ_MODE0 = 1'b0;
defparam dpx9b_inst_18.READ_MODE1 = 1'b0;
defparam dpx9b_inst_18.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_18.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_18.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_18.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_18.BLK_SEL_0 = 3'b010;
defparam dpx9b_inst_18.BLK_SEL_1 = 3'b010;
defparam dpx9b_inst_18.RESET_MODE = "SYNC";
defparam dpx9b_inst_18.INIT_RAM_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_18.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_19 (
    .DOA({dpx9b_inst_19_douta_w[8:0],dpx9b_inst_19_douta[26:18]}),
    .DOB({dpx9b_inst_19_doutb_w[8:0],dpx9b_inst_19_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_19.READ_MODE0 = 1'b0;
defparam dpx9b_inst_19.READ_MODE1 = 1'b0;
defparam dpx9b_inst_19.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_19.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_19.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_19.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_19.BLK_SEL_0 = 3'b011;
defparam dpx9b_inst_19.BLK_SEL_1 = 3'b011;
defparam dpx9b_inst_19.RESET_MODE = "SYNC";
defparam dpx9b_inst_19.INIT_RAM_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_19.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_20 (
    .DOA({dpx9b_inst_20_douta_w[8:0],dpx9b_inst_20_douta[26:18]}),
    .DOB({dpx9b_inst_20_doutb_w[8:0],dpx9b_inst_20_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_20.READ_MODE0 = 1'b0;
defparam dpx9b_inst_20.READ_MODE1 = 1'b0;
defparam dpx9b_inst_20.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_20.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_20.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_20.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_20.BLK_SEL_0 = 3'b100;
defparam dpx9b_inst_20.BLK_SEL_1 = 3'b100;
defparam dpx9b_inst_20.RESET_MODE = "SYNC";
defparam dpx9b_inst_20.INIT_RAM_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_20.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_21 (
    .DOA({dpx9b_inst_21_douta_w[8:0],dpx9b_inst_21_douta[26:18]}),
    .DOB({dpx9b_inst_21_doutb_w[8:0],dpx9b_inst_21_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_21.READ_MODE0 = 1'b0;
defparam dpx9b_inst_21.READ_MODE1 = 1'b0;
defparam dpx9b_inst_21.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_21.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_21.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_21.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_21.BLK_SEL_0 = 3'b101;
defparam dpx9b_inst_21.BLK_SEL_1 = 3'b101;
defparam dpx9b_inst_21.RESET_MODE = "SYNC";
defparam dpx9b_inst_21.INIT_RAM_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_21.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_22 (
    .DOA({dpx9b_inst_22_douta_w[8:0],dpx9b_inst_22_douta[26:18]}),
    .DOB({dpx9b_inst_22_doutb_w[8:0],dpx9b_inst_22_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_22.READ_MODE0 = 1'b0;
defparam dpx9b_inst_22.READ_MODE1 = 1'b0;
defparam dpx9b_inst_22.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_22.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_22.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_22.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_22.BLK_SEL_0 = 3'b110;
defparam dpx9b_inst_22.BLK_SEL_1 = 3'b110;
defparam dpx9b_inst_22.RESET_MODE = "SYNC";
defparam dpx9b_inst_22.INIT_RAM_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_22.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPX9B dpx9b_inst_23 (
    .DOA({dpx9b_inst_23_douta_w[8:0],dpx9b_inst_23_douta[26:18]}),
    .DOB({dpx9b_inst_23_doutb_w[8:0],dpx9b_inst_23_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_23.READ_MODE0 = 1'b0;
defparam dpx9b_inst_23.READ_MODE1 = 1'b0;
defparam dpx9b_inst_23.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_23.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_23.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_23.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_23.BLK_SEL_0 = 3'b111;
defparam dpx9b_inst_23.BLK_SEL_1 = 3'b111;
defparam dpx9b_inst_23.RESET_MODE = "SYNC";
defparam dpx9b_inst_23.INIT_RAM_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam dpx9b_inst_23.INIT_RAM_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_24 (
    .DOA({dpb_inst_24_douta_w[14:0],douta[27]}),
    .DOB({dpb_inst_24_doutb_w[14:0],doutb[27]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[27]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[27]})
);

defparam dpb_inst_24.READ_MODE0 = 1'b0;
defparam dpb_inst_24.READ_MODE1 = 1'b0;
defparam dpb_inst_24.WRITE_MODE0 = 2'b00;
defparam dpb_inst_24.WRITE_MODE1 = 2'b00;
defparam dpb_inst_24.BIT_WIDTH_0 = 1;
defparam dpb_inst_24.BIT_WIDTH_1 = 1;
defparam dpb_inst_24.BLK_SEL_0 = 3'b000;
defparam dpb_inst_24.BLK_SEL_1 = 3'b000;
defparam dpb_inst_24.RESET_MODE = "SYNC";
defparam dpb_inst_24.INIT_RAM_00 = 256'h5810080891A5462C0888605E9D120448D0216C818C656260800000002DA18800;
defparam dpb_inst_24.INIT_RAM_01 = 256'h0000000000001FFFFFFFE00000000043434308530A85080808C0808D0A3468D6;
defparam dpb_inst_24.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_0B = 256'h0200C4C080000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_0C = 256'h000000000000000000000000000000000000000000000000062C480224880312;
defparam dpb_inst_24.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_24.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_25 (
    .DOA({dpb_inst_25_douta_w[14:0],douta[28]}),
    .DOB({dpb_inst_25_doutb_w[14:0],doutb[28]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[28]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[28]})
);

defparam dpb_inst_25.READ_MODE0 = 1'b0;
defparam dpb_inst_25.READ_MODE1 = 1'b0;
defparam dpb_inst_25.WRITE_MODE0 = 2'b00;
defparam dpb_inst_25.WRITE_MODE1 = 2'b00;
defparam dpb_inst_25.BIT_WIDTH_0 = 1;
defparam dpb_inst_25.BIT_WIDTH_1 = 1;
defparam dpb_inst_25.BLK_SEL_0 = 3'b000;
defparam dpb_inst_25.BLK_SEL_1 = 3'b000;
defparam dpb_inst_25.RESET_MODE = "SYNC";
defparam dpb_inst_25.INIT_RAM_00 = 256'h810D348040040440804AC41A140840200201421000020C0F01AD1BA0508A8040;
defparam dpb_inst_25.INIT_RAM_01 = 256'h000000000000000000000000000003151515020D052C9134805B480400102048;
defparam dpb_inst_25.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_0B = 256'hD200F8F480000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_0C = 256'h00000000000000000000000000000000000000000000000007CFA803C76803E3;
defparam dpb_inst_25.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_25.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_26 (
    .DOA({dpb_inst_26_douta_w[14:0],douta[29]}),
    .DOB({dpb_inst_26_doutb_w[14:0],doutb[29]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[29]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[29]})
);

defparam dpb_inst_26.READ_MODE0 = 1'b0;
defparam dpb_inst_26.READ_MODE1 = 1'b0;
defparam dpb_inst_26.WRITE_MODE0 = 2'b00;
defparam dpb_inst_26.WRITE_MODE1 = 2'b00;
defparam dpb_inst_26.BIT_WIDTH_0 = 1;
defparam dpb_inst_26.BIT_WIDTH_1 = 1;
defparam dpb_inst_26.BLK_SEL_0 = 3'b000;
defparam dpb_inst_26.BLK_SEL_1 = 3'b000;
defparam dpb_inst_26.RESET_MODE = "SYNC";
defparam dpb_inst_26.INIT_RAM_00 = 256'hFFDC43E7CF9D3EFFE7D33F2C78F9F3E7CF9E7FFDDEF3FF7FFDFFDFFBFF903DEC;
defparam dpb_inst_26.INIT_RAM_01 = 256'h00000000000000000000000000000330303074B37CBFB443E7843E78F9E3C79F;
defparam dpb_inst_26.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_0B = 256'h0200000080000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000280000280000;
defparam dpb_inst_26.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_26.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_27 (
    .DOA({dpb_inst_27_douta_w[14:0],douta[30]}),
    .DOB({dpb_inst_27_doutb_w[14:0],doutb[30]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[30]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[30]})
);

defparam dpb_inst_27.READ_MODE0 = 1'b0;
defparam dpb_inst_27.READ_MODE1 = 1'b0;
defparam dpb_inst_27.WRITE_MODE0 = 2'b00;
defparam dpb_inst_27.WRITE_MODE1 = 2'b00;
defparam dpb_inst_27.BIT_WIDTH_0 = 1;
defparam dpb_inst_27.BIT_WIDTH_1 = 1;
defparam dpb_inst_27.BLK_SEL_0 = 3'b000;
defparam dpb_inst_27.BLK_SEL_1 = 3'b000;
defparam dpb_inst_27.RESET_MODE = "SYNC";
defparam dpb_inst_27.INIT_RAM_00 = 256'hFB1DBD80C18302FD80D8EC160C10C040C6033F9DCC63FF7FCDBF5BE9B7AFA940;
defparam dpb_inst_27.INIT_RAM_01 = 256'h00000000000000000000000000000C4F4F4F6E7F0FBD9DBD80DBD80C183060DD;
defparam dpb_inst_27.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_0B = 256'h0A01FE0280000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000FE00807F00807F8;
defparam dpb_inst_27.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_27.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_28 (
    .DOA({dpb_inst_28_douta_w[14:0],douta[31]}),
    .DOB({dpb_inst_28_doutb_w[14:0],doutb[31]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[31]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[31]})
);

defparam dpb_inst_28.READ_MODE0 = 1'b0;
defparam dpb_inst_28.READ_MODE1 = 1'b0;
defparam dpb_inst_28.WRITE_MODE0 = 2'b00;
defparam dpb_inst_28.WRITE_MODE1 = 2'b00;
defparam dpb_inst_28.BIT_WIDTH_0 = 1;
defparam dpb_inst_28.BIT_WIDTH_1 = 1;
defparam dpb_inst_28.BLK_SEL_0 = 3'b000;
defparam dpb_inst_28.BLK_SEL_1 = 3'b000;
defparam dpb_inst_28.RESET_MODE = "SYNC";
defparam dpb_inst_28.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_0B = 256'hF200FEFC80000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_0C = 256'h00000000000000000000000000000000000000000000000007EFC803F7C803FB;
defparam dpb_inst_28.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_28.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ada[13]),
  .CLK(clka),
  .CE(cea_w)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(ada[12]),
  .CLK(clka),
  .CE(cea_w)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(ada[11]),
  .CLK(clka),
  .CE(cea_w)
);
DFFE dff_inst_3 (
  .Q(dff_q_3),
  .D(adb[13]),
  .CLK(clkb),
  .CE(ceb_w)
);
DFFE dff_inst_4 (
  .Q(dff_q_4),
  .D(adb[12]),
  .CLK(clkb),
  .CE(ceb_w)
);
DFFE dff_inst_5 (
  .Q(dff_q_5),
  .D(adb[11]),
  .CLK(clkb),
  .CE(ceb_w)
);
MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(dpx9b_inst_0_douta[0]),
  .I1(dpx9b_inst_1_douta[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(dpx9b_inst_2_douta[0]),
  .I1(dpx9b_inst_3_douta[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(dpx9b_inst_4_douta[0]),
  .I1(dpx9b_inst_5_douta[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(dpx9b_inst_6_douta[0]),
  .I1(dpx9b_inst_7_douta[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(dff_q_1)
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(dff_q_1)
);
MUX2 mux_inst_6 (
  .O(douta[0]),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(dff_q_0)
);
MUX2 mux_inst_7 (
  .O(mux_o_7),
  .I0(dpx9b_inst_0_douta[1]),
  .I1(dpx9b_inst_1_douta[1]),
  .S0(dff_q_2)
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(dpx9b_inst_2_douta[1]),
  .I1(dpx9b_inst_3_douta[1]),
  .S0(dff_q_2)
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(dpx9b_inst_4_douta[1]),
  .I1(dpx9b_inst_5_douta[1]),
  .S0(dff_q_2)
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(dpx9b_inst_6_douta[1]),
  .I1(dpx9b_inst_7_douta[1]),
  .S0(dff_q_2)
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(mux_o_7),
  .I1(mux_o_8),
  .S0(dff_q_1)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(mux_o_9),
  .I1(mux_o_10),
  .S0(dff_q_1)
);
MUX2 mux_inst_13 (
  .O(douta[1]),
  .I0(mux_o_11),
  .I1(mux_o_12),
  .S0(dff_q_0)
);
MUX2 mux_inst_14 (
  .O(mux_o_14),
  .I0(dpx9b_inst_0_douta[2]),
  .I1(dpx9b_inst_1_douta[2]),
  .S0(dff_q_2)
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(dpx9b_inst_2_douta[2]),
  .I1(dpx9b_inst_3_douta[2]),
  .S0(dff_q_2)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(dpx9b_inst_4_douta[2]),
  .I1(dpx9b_inst_5_douta[2]),
  .S0(dff_q_2)
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(dpx9b_inst_6_douta[2]),
  .I1(dpx9b_inst_7_douta[2]),
  .S0(dff_q_2)
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(mux_o_14),
  .I1(mux_o_15),
  .S0(dff_q_1)
);
MUX2 mux_inst_19 (
  .O(mux_o_19),
  .I0(mux_o_16),
  .I1(mux_o_17),
  .S0(dff_q_1)
);
MUX2 mux_inst_20 (
  .O(douta[2]),
  .I0(mux_o_18),
  .I1(mux_o_19),
  .S0(dff_q_0)
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(dpx9b_inst_0_douta[3]),
  .I1(dpx9b_inst_1_douta[3]),
  .S0(dff_q_2)
);
MUX2 mux_inst_22 (
  .O(mux_o_22),
  .I0(dpx9b_inst_2_douta[3]),
  .I1(dpx9b_inst_3_douta[3]),
  .S0(dff_q_2)
);
MUX2 mux_inst_23 (
  .O(mux_o_23),
  .I0(dpx9b_inst_4_douta[3]),
  .I1(dpx9b_inst_5_douta[3]),
  .S0(dff_q_2)
);
MUX2 mux_inst_24 (
  .O(mux_o_24),
  .I0(dpx9b_inst_6_douta[3]),
  .I1(dpx9b_inst_7_douta[3]),
  .S0(dff_q_2)
);
MUX2 mux_inst_25 (
  .O(mux_o_25),
  .I0(mux_o_21),
  .I1(mux_o_22),
  .S0(dff_q_1)
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(mux_o_23),
  .I1(mux_o_24),
  .S0(dff_q_1)
);
MUX2 mux_inst_27 (
  .O(douta[3]),
  .I0(mux_o_25),
  .I1(mux_o_26),
  .S0(dff_q_0)
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(dpx9b_inst_0_douta[4]),
  .I1(dpx9b_inst_1_douta[4]),
  .S0(dff_q_2)
);
MUX2 mux_inst_29 (
  .O(mux_o_29),
  .I0(dpx9b_inst_2_douta[4]),
  .I1(dpx9b_inst_3_douta[4]),
  .S0(dff_q_2)
);
MUX2 mux_inst_30 (
  .O(mux_o_30),
  .I0(dpx9b_inst_4_douta[4]),
  .I1(dpx9b_inst_5_douta[4]),
  .S0(dff_q_2)
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(dpx9b_inst_6_douta[4]),
  .I1(dpx9b_inst_7_douta[4]),
  .S0(dff_q_2)
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(mux_o_28),
  .I1(mux_o_29),
  .S0(dff_q_1)
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(mux_o_30),
  .I1(mux_o_31),
  .S0(dff_q_1)
);
MUX2 mux_inst_34 (
  .O(douta[4]),
  .I0(mux_o_32),
  .I1(mux_o_33),
  .S0(dff_q_0)
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(dpx9b_inst_0_douta[5]),
  .I1(dpx9b_inst_1_douta[5]),
  .S0(dff_q_2)
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(dpx9b_inst_2_douta[5]),
  .I1(dpx9b_inst_3_douta[5]),
  .S0(dff_q_2)
);
MUX2 mux_inst_37 (
  .O(mux_o_37),
  .I0(dpx9b_inst_4_douta[5]),
  .I1(dpx9b_inst_5_douta[5]),
  .S0(dff_q_2)
);
MUX2 mux_inst_38 (
  .O(mux_o_38),
  .I0(dpx9b_inst_6_douta[5]),
  .I1(dpx9b_inst_7_douta[5]),
  .S0(dff_q_2)
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(mux_o_35),
  .I1(mux_o_36),
  .S0(dff_q_1)
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(mux_o_37),
  .I1(mux_o_38),
  .S0(dff_q_1)
);
MUX2 mux_inst_41 (
  .O(douta[5]),
  .I0(mux_o_39),
  .I1(mux_o_40),
  .S0(dff_q_0)
);
MUX2 mux_inst_42 (
  .O(mux_o_42),
  .I0(dpx9b_inst_0_douta[6]),
  .I1(dpx9b_inst_1_douta[6]),
  .S0(dff_q_2)
);
MUX2 mux_inst_43 (
  .O(mux_o_43),
  .I0(dpx9b_inst_2_douta[6]),
  .I1(dpx9b_inst_3_douta[6]),
  .S0(dff_q_2)
);
MUX2 mux_inst_44 (
  .O(mux_o_44),
  .I0(dpx9b_inst_4_douta[6]),
  .I1(dpx9b_inst_5_douta[6]),
  .S0(dff_q_2)
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(dpx9b_inst_6_douta[6]),
  .I1(dpx9b_inst_7_douta[6]),
  .S0(dff_q_2)
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(mux_o_42),
  .I1(mux_o_43),
  .S0(dff_q_1)
);
MUX2 mux_inst_47 (
  .O(mux_o_47),
  .I0(mux_o_44),
  .I1(mux_o_45),
  .S0(dff_q_1)
);
MUX2 mux_inst_48 (
  .O(douta[6]),
  .I0(mux_o_46),
  .I1(mux_o_47),
  .S0(dff_q_0)
);
MUX2 mux_inst_49 (
  .O(mux_o_49),
  .I0(dpx9b_inst_0_douta[7]),
  .I1(dpx9b_inst_1_douta[7]),
  .S0(dff_q_2)
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(dpx9b_inst_2_douta[7]),
  .I1(dpx9b_inst_3_douta[7]),
  .S0(dff_q_2)
);
MUX2 mux_inst_51 (
  .O(mux_o_51),
  .I0(dpx9b_inst_4_douta[7]),
  .I1(dpx9b_inst_5_douta[7]),
  .S0(dff_q_2)
);
MUX2 mux_inst_52 (
  .O(mux_o_52),
  .I0(dpx9b_inst_6_douta[7]),
  .I1(dpx9b_inst_7_douta[7]),
  .S0(dff_q_2)
);
MUX2 mux_inst_53 (
  .O(mux_o_53),
  .I0(mux_o_49),
  .I1(mux_o_50),
  .S0(dff_q_1)
);
MUX2 mux_inst_54 (
  .O(mux_o_54),
  .I0(mux_o_51),
  .I1(mux_o_52),
  .S0(dff_q_1)
);
MUX2 mux_inst_55 (
  .O(douta[7]),
  .I0(mux_o_53),
  .I1(mux_o_54),
  .S0(dff_q_0)
);
MUX2 mux_inst_56 (
  .O(mux_o_56),
  .I0(dpx9b_inst_0_douta[8]),
  .I1(dpx9b_inst_1_douta[8]),
  .S0(dff_q_2)
);
MUX2 mux_inst_57 (
  .O(mux_o_57),
  .I0(dpx9b_inst_2_douta[8]),
  .I1(dpx9b_inst_3_douta[8]),
  .S0(dff_q_2)
);
MUX2 mux_inst_58 (
  .O(mux_o_58),
  .I0(dpx9b_inst_4_douta[8]),
  .I1(dpx9b_inst_5_douta[8]),
  .S0(dff_q_2)
);
MUX2 mux_inst_59 (
  .O(mux_o_59),
  .I0(dpx9b_inst_6_douta[8]),
  .I1(dpx9b_inst_7_douta[8]),
  .S0(dff_q_2)
);
MUX2 mux_inst_60 (
  .O(mux_o_60),
  .I0(mux_o_56),
  .I1(mux_o_57),
  .S0(dff_q_1)
);
MUX2 mux_inst_61 (
  .O(mux_o_61),
  .I0(mux_o_58),
  .I1(mux_o_59),
  .S0(dff_q_1)
);
MUX2 mux_inst_62 (
  .O(douta[8]),
  .I0(mux_o_60),
  .I1(mux_o_61),
  .S0(dff_q_0)
);
MUX2 mux_inst_63 (
  .O(mux_o_63),
  .I0(dpx9b_inst_8_douta[9]),
  .I1(dpx9b_inst_9_douta[9]),
  .S0(dff_q_2)
);
MUX2 mux_inst_64 (
  .O(mux_o_64),
  .I0(dpx9b_inst_10_douta[9]),
  .I1(dpx9b_inst_11_douta[9]),
  .S0(dff_q_2)
);
MUX2 mux_inst_65 (
  .O(mux_o_65),
  .I0(dpx9b_inst_12_douta[9]),
  .I1(dpx9b_inst_13_douta[9]),
  .S0(dff_q_2)
);
MUX2 mux_inst_66 (
  .O(mux_o_66),
  .I0(dpx9b_inst_14_douta[9]),
  .I1(dpx9b_inst_15_douta[9]),
  .S0(dff_q_2)
);
MUX2 mux_inst_67 (
  .O(mux_o_67),
  .I0(mux_o_63),
  .I1(mux_o_64),
  .S0(dff_q_1)
);
MUX2 mux_inst_68 (
  .O(mux_o_68),
  .I0(mux_o_65),
  .I1(mux_o_66),
  .S0(dff_q_1)
);
MUX2 mux_inst_69 (
  .O(douta[9]),
  .I0(mux_o_67),
  .I1(mux_o_68),
  .S0(dff_q_0)
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(dpx9b_inst_8_douta[10]),
  .I1(dpx9b_inst_9_douta[10]),
  .S0(dff_q_2)
);
MUX2 mux_inst_71 (
  .O(mux_o_71),
  .I0(dpx9b_inst_10_douta[10]),
  .I1(dpx9b_inst_11_douta[10]),
  .S0(dff_q_2)
);
MUX2 mux_inst_72 (
  .O(mux_o_72),
  .I0(dpx9b_inst_12_douta[10]),
  .I1(dpx9b_inst_13_douta[10]),
  .S0(dff_q_2)
);
MUX2 mux_inst_73 (
  .O(mux_o_73),
  .I0(dpx9b_inst_14_douta[10]),
  .I1(dpx9b_inst_15_douta[10]),
  .S0(dff_q_2)
);
MUX2 mux_inst_74 (
  .O(mux_o_74),
  .I0(mux_o_70),
  .I1(mux_o_71),
  .S0(dff_q_1)
);
MUX2 mux_inst_75 (
  .O(mux_o_75),
  .I0(mux_o_72),
  .I1(mux_o_73),
  .S0(dff_q_1)
);
MUX2 mux_inst_76 (
  .O(douta[10]),
  .I0(mux_o_74),
  .I1(mux_o_75),
  .S0(dff_q_0)
);
MUX2 mux_inst_77 (
  .O(mux_o_77),
  .I0(dpx9b_inst_8_douta[11]),
  .I1(dpx9b_inst_9_douta[11]),
  .S0(dff_q_2)
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(dpx9b_inst_10_douta[11]),
  .I1(dpx9b_inst_11_douta[11]),
  .S0(dff_q_2)
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(dpx9b_inst_12_douta[11]),
  .I1(dpx9b_inst_13_douta[11]),
  .S0(dff_q_2)
);
MUX2 mux_inst_80 (
  .O(mux_o_80),
  .I0(dpx9b_inst_14_douta[11]),
  .I1(dpx9b_inst_15_douta[11]),
  .S0(dff_q_2)
);
MUX2 mux_inst_81 (
  .O(mux_o_81),
  .I0(mux_o_77),
  .I1(mux_o_78),
  .S0(dff_q_1)
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(mux_o_79),
  .I1(mux_o_80),
  .S0(dff_q_1)
);
MUX2 mux_inst_83 (
  .O(douta[11]),
  .I0(mux_o_81),
  .I1(mux_o_82),
  .S0(dff_q_0)
);
MUX2 mux_inst_84 (
  .O(mux_o_84),
  .I0(dpx9b_inst_8_douta[12]),
  .I1(dpx9b_inst_9_douta[12]),
  .S0(dff_q_2)
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(dpx9b_inst_10_douta[12]),
  .I1(dpx9b_inst_11_douta[12]),
  .S0(dff_q_2)
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(dpx9b_inst_12_douta[12]),
  .I1(dpx9b_inst_13_douta[12]),
  .S0(dff_q_2)
);
MUX2 mux_inst_87 (
  .O(mux_o_87),
  .I0(dpx9b_inst_14_douta[12]),
  .I1(dpx9b_inst_15_douta[12]),
  .S0(dff_q_2)
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(mux_o_84),
  .I1(mux_o_85),
  .S0(dff_q_1)
);
MUX2 mux_inst_89 (
  .O(mux_o_89),
  .I0(mux_o_86),
  .I1(mux_o_87),
  .S0(dff_q_1)
);
MUX2 mux_inst_90 (
  .O(douta[12]),
  .I0(mux_o_88),
  .I1(mux_o_89),
  .S0(dff_q_0)
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(dpx9b_inst_8_douta[13]),
  .I1(dpx9b_inst_9_douta[13]),
  .S0(dff_q_2)
);
MUX2 mux_inst_92 (
  .O(mux_o_92),
  .I0(dpx9b_inst_10_douta[13]),
  .I1(dpx9b_inst_11_douta[13]),
  .S0(dff_q_2)
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(dpx9b_inst_12_douta[13]),
  .I1(dpx9b_inst_13_douta[13]),
  .S0(dff_q_2)
);
MUX2 mux_inst_94 (
  .O(mux_o_94),
  .I0(dpx9b_inst_14_douta[13]),
  .I1(dpx9b_inst_15_douta[13]),
  .S0(dff_q_2)
);
MUX2 mux_inst_95 (
  .O(mux_o_95),
  .I0(mux_o_91),
  .I1(mux_o_92),
  .S0(dff_q_1)
);
MUX2 mux_inst_96 (
  .O(mux_o_96),
  .I0(mux_o_93),
  .I1(mux_o_94),
  .S0(dff_q_1)
);
MUX2 mux_inst_97 (
  .O(douta[13]),
  .I0(mux_o_95),
  .I1(mux_o_96),
  .S0(dff_q_0)
);
MUX2 mux_inst_98 (
  .O(mux_o_98),
  .I0(dpx9b_inst_8_douta[14]),
  .I1(dpx9b_inst_9_douta[14]),
  .S0(dff_q_2)
);
MUX2 mux_inst_99 (
  .O(mux_o_99),
  .I0(dpx9b_inst_10_douta[14]),
  .I1(dpx9b_inst_11_douta[14]),
  .S0(dff_q_2)
);
MUX2 mux_inst_100 (
  .O(mux_o_100),
  .I0(dpx9b_inst_12_douta[14]),
  .I1(dpx9b_inst_13_douta[14]),
  .S0(dff_q_2)
);
MUX2 mux_inst_101 (
  .O(mux_o_101),
  .I0(dpx9b_inst_14_douta[14]),
  .I1(dpx9b_inst_15_douta[14]),
  .S0(dff_q_2)
);
MUX2 mux_inst_102 (
  .O(mux_o_102),
  .I0(mux_o_98),
  .I1(mux_o_99),
  .S0(dff_q_1)
);
MUX2 mux_inst_103 (
  .O(mux_o_103),
  .I0(mux_o_100),
  .I1(mux_o_101),
  .S0(dff_q_1)
);
MUX2 mux_inst_104 (
  .O(douta[14]),
  .I0(mux_o_102),
  .I1(mux_o_103),
  .S0(dff_q_0)
);
MUX2 mux_inst_105 (
  .O(mux_o_105),
  .I0(dpx9b_inst_8_douta[15]),
  .I1(dpx9b_inst_9_douta[15]),
  .S0(dff_q_2)
);
MUX2 mux_inst_106 (
  .O(mux_o_106),
  .I0(dpx9b_inst_10_douta[15]),
  .I1(dpx9b_inst_11_douta[15]),
  .S0(dff_q_2)
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(dpx9b_inst_12_douta[15]),
  .I1(dpx9b_inst_13_douta[15]),
  .S0(dff_q_2)
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(dpx9b_inst_14_douta[15]),
  .I1(dpx9b_inst_15_douta[15]),
  .S0(dff_q_2)
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(mux_o_105),
  .I1(mux_o_106),
  .S0(dff_q_1)
);
MUX2 mux_inst_110 (
  .O(mux_o_110),
  .I0(mux_o_107),
  .I1(mux_o_108),
  .S0(dff_q_1)
);
MUX2 mux_inst_111 (
  .O(douta[15]),
  .I0(mux_o_109),
  .I1(mux_o_110),
  .S0(dff_q_0)
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(dpx9b_inst_8_douta[16]),
  .I1(dpx9b_inst_9_douta[16]),
  .S0(dff_q_2)
);
MUX2 mux_inst_113 (
  .O(mux_o_113),
  .I0(dpx9b_inst_10_douta[16]),
  .I1(dpx9b_inst_11_douta[16]),
  .S0(dff_q_2)
);
MUX2 mux_inst_114 (
  .O(mux_o_114),
  .I0(dpx9b_inst_12_douta[16]),
  .I1(dpx9b_inst_13_douta[16]),
  .S0(dff_q_2)
);
MUX2 mux_inst_115 (
  .O(mux_o_115),
  .I0(dpx9b_inst_14_douta[16]),
  .I1(dpx9b_inst_15_douta[16]),
  .S0(dff_q_2)
);
MUX2 mux_inst_116 (
  .O(mux_o_116),
  .I0(mux_o_112),
  .I1(mux_o_113),
  .S0(dff_q_1)
);
MUX2 mux_inst_117 (
  .O(mux_o_117),
  .I0(mux_o_114),
  .I1(mux_o_115),
  .S0(dff_q_1)
);
MUX2 mux_inst_118 (
  .O(douta[16]),
  .I0(mux_o_116),
  .I1(mux_o_117),
  .S0(dff_q_0)
);
MUX2 mux_inst_119 (
  .O(mux_o_119),
  .I0(dpx9b_inst_8_douta[17]),
  .I1(dpx9b_inst_9_douta[17]),
  .S0(dff_q_2)
);
MUX2 mux_inst_120 (
  .O(mux_o_120),
  .I0(dpx9b_inst_10_douta[17]),
  .I1(dpx9b_inst_11_douta[17]),
  .S0(dff_q_2)
);
MUX2 mux_inst_121 (
  .O(mux_o_121),
  .I0(dpx9b_inst_12_douta[17]),
  .I1(dpx9b_inst_13_douta[17]),
  .S0(dff_q_2)
);
MUX2 mux_inst_122 (
  .O(mux_o_122),
  .I0(dpx9b_inst_14_douta[17]),
  .I1(dpx9b_inst_15_douta[17]),
  .S0(dff_q_2)
);
MUX2 mux_inst_123 (
  .O(mux_o_123),
  .I0(mux_o_119),
  .I1(mux_o_120),
  .S0(dff_q_1)
);
MUX2 mux_inst_124 (
  .O(mux_o_124),
  .I0(mux_o_121),
  .I1(mux_o_122),
  .S0(dff_q_1)
);
MUX2 mux_inst_125 (
  .O(douta[17]),
  .I0(mux_o_123),
  .I1(mux_o_124),
  .S0(dff_q_0)
);
MUX2 mux_inst_126 (
  .O(mux_o_126),
  .I0(dpx9b_inst_16_douta[18]),
  .I1(dpx9b_inst_17_douta[18]),
  .S0(dff_q_2)
);
MUX2 mux_inst_127 (
  .O(mux_o_127),
  .I0(dpx9b_inst_18_douta[18]),
  .I1(dpx9b_inst_19_douta[18]),
  .S0(dff_q_2)
);
MUX2 mux_inst_128 (
  .O(mux_o_128),
  .I0(dpx9b_inst_20_douta[18]),
  .I1(dpx9b_inst_21_douta[18]),
  .S0(dff_q_2)
);
MUX2 mux_inst_129 (
  .O(mux_o_129),
  .I0(dpx9b_inst_22_douta[18]),
  .I1(dpx9b_inst_23_douta[18]),
  .S0(dff_q_2)
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(mux_o_126),
  .I1(mux_o_127),
  .S0(dff_q_1)
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(mux_o_128),
  .I1(mux_o_129),
  .S0(dff_q_1)
);
MUX2 mux_inst_132 (
  .O(douta[18]),
  .I0(mux_o_130),
  .I1(mux_o_131),
  .S0(dff_q_0)
);
MUX2 mux_inst_133 (
  .O(mux_o_133),
  .I0(dpx9b_inst_16_douta[19]),
  .I1(dpx9b_inst_17_douta[19]),
  .S0(dff_q_2)
);
MUX2 mux_inst_134 (
  .O(mux_o_134),
  .I0(dpx9b_inst_18_douta[19]),
  .I1(dpx9b_inst_19_douta[19]),
  .S0(dff_q_2)
);
MUX2 mux_inst_135 (
  .O(mux_o_135),
  .I0(dpx9b_inst_20_douta[19]),
  .I1(dpx9b_inst_21_douta[19]),
  .S0(dff_q_2)
);
MUX2 mux_inst_136 (
  .O(mux_o_136),
  .I0(dpx9b_inst_22_douta[19]),
  .I1(dpx9b_inst_23_douta[19]),
  .S0(dff_q_2)
);
MUX2 mux_inst_137 (
  .O(mux_o_137),
  .I0(mux_o_133),
  .I1(mux_o_134),
  .S0(dff_q_1)
);
MUX2 mux_inst_138 (
  .O(mux_o_138),
  .I0(mux_o_135),
  .I1(mux_o_136),
  .S0(dff_q_1)
);
MUX2 mux_inst_139 (
  .O(douta[19]),
  .I0(mux_o_137),
  .I1(mux_o_138),
  .S0(dff_q_0)
);
MUX2 mux_inst_140 (
  .O(mux_o_140),
  .I0(dpx9b_inst_16_douta[20]),
  .I1(dpx9b_inst_17_douta[20]),
  .S0(dff_q_2)
);
MUX2 mux_inst_141 (
  .O(mux_o_141),
  .I0(dpx9b_inst_18_douta[20]),
  .I1(dpx9b_inst_19_douta[20]),
  .S0(dff_q_2)
);
MUX2 mux_inst_142 (
  .O(mux_o_142),
  .I0(dpx9b_inst_20_douta[20]),
  .I1(dpx9b_inst_21_douta[20]),
  .S0(dff_q_2)
);
MUX2 mux_inst_143 (
  .O(mux_o_143),
  .I0(dpx9b_inst_22_douta[20]),
  .I1(dpx9b_inst_23_douta[20]),
  .S0(dff_q_2)
);
MUX2 mux_inst_144 (
  .O(mux_o_144),
  .I0(mux_o_140),
  .I1(mux_o_141),
  .S0(dff_q_1)
);
MUX2 mux_inst_145 (
  .O(mux_o_145),
  .I0(mux_o_142),
  .I1(mux_o_143),
  .S0(dff_q_1)
);
MUX2 mux_inst_146 (
  .O(douta[20]),
  .I0(mux_o_144),
  .I1(mux_o_145),
  .S0(dff_q_0)
);
MUX2 mux_inst_147 (
  .O(mux_o_147),
  .I0(dpx9b_inst_16_douta[21]),
  .I1(dpx9b_inst_17_douta[21]),
  .S0(dff_q_2)
);
MUX2 mux_inst_148 (
  .O(mux_o_148),
  .I0(dpx9b_inst_18_douta[21]),
  .I1(dpx9b_inst_19_douta[21]),
  .S0(dff_q_2)
);
MUX2 mux_inst_149 (
  .O(mux_o_149),
  .I0(dpx9b_inst_20_douta[21]),
  .I1(dpx9b_inst_21_douta[21]),
  .S0(dff_q_2)
);
MUX2 mux_inst_150 (
  .O(mux_o_150),
  .I0(dpx9b_inst_22_douta[21]),
  .I1(dpx9b_inst_23_douta[21]),
  .S0(dff_q_2)
);
MUX2 mux_inst_151 (
  .O(mux_o_151),
  .I0(mux_o_147),
  .I1(mux_o_148),
  .S0(dff_q_1)
);
MUX2 mux_inst_152 (
  .O(mux_o_152),
  .I0(mux_o_149),
  .I1(mux_o_150),
  .S0(dff_q_1)
);
MUX2 mux_inst_153 (
  .O(douta[21]),
  .I0(mux_o_151),
  .I1(mux_o_152),
  .S0(dff_q_0)
);
MUX2 mux_inst_154 (
  .O(mux_o_154),
  .I0(dpx9b_inst_16_douta[22]),
  .I1(dpx9b_inst_17_douta[22]),
  .S0(dff_q_2)
);
MUX2 mux_inst_155 (
  .O(mux_o_155),
  .I0(dpx9b_inst_18_douta[22]),
  .I1(dpx9b_inst_19_douta[22]),
  .S0(dff_q_2)
);
MUX2 mux_inst_156 (
  .O(mux_o_156),
  .I0(dpx9b_inst_20_douta[22]),
  .I1(dpx9b_inst_21_douta[22]),
  .S0(dff_q_2)
);
MUX2 mux_inst_157 (
  .O(mux_o_157),
  .I0(dpx9b_inst_22_douta[22]),
  .I1(dpx9b_inst_23_douta[22]),
  .S0(dff_q_2)
);
MUX2 mux_inst_158 (
  .O(mux_o_158),
  .I0(mux_o_154),
  .I1(mux_o_155),
  .S0(dff_q_1)
);
MUX2 mux_inst_159 (
  .O(mux_o_159),
  .I0(mux_o_156),
  .I1(mux_o_157),
  .S0(dff_q_1)
);
MUX2 mux_inst_160 (
  .O(douta[22]),
  .I0(mux_o_158),
  .I1(mux_o_159),
  .S0(dff_q_0)
);
MUX2 mux_inst_161 (
  .O(mux_o_161),
  .I0(dpx9b_inst_16_douta[23]),
  .I1(dpx9b_inst_17_douta[23]),
  .S0(dff_q_2)
);
MUX2 mux_inst_162 (
  .O(mux_o_162),
  .I0(dpx9b_inst_18_douta[23]),
  .I1(dpx9b_inst_19_douta[23]),
  .S0(dff_q_2)
);
MUX2 mux_inst_163 (
  .O(mux_o_163),
  .I0(dpx9b_inst_20_douta[23]),
  .I1(dpx9b_inst_21_douta[23]),
  .S0(dff_q_2)
);
MUX2 mux_inst_164 (
  .O(mux_o_164),
  .I0(dpx9b_inst_22_douta[23]),
  .I1(dpx9b_inst_23_douta[23]),
  .S0(dff_q_2)
);
MUX2 mux_inst_165 (
  .O(mux_o_165),
  .I0(mux_o_161),
  .I1(mux_o_162),
  .S0(dff_q_1)
);
MUX2 mux_inst_166 (
  .O(mux_o_166),
  .I0(mux_o_163),
  .I1(mux_o_164),
  .S0(dff_q_1)
);
MUX2 mux_inst_167 (
  .O(douta[23]),
  .I0(mux_o_165),
  .I1(mux_o_166),
  .S0(dff_q_0)
);
MUX2 mux_inst_168 (
  .O(mux_o_168),
  .I0(dpx9b_inst_16_douta[24]),
  .I1(dpx9b_inst_17_douta[24]),
  .S0(dff_q_2)
);
MUX2 mux_inst_169 (
  .O(mux_o_169),
  .I0(dpx9b_inst_18_douta[24]),
  .I1(dpx9b_inst_19_douta[24]),
  .S0(dff_q_2)
);
MUX2 mux_inst_170 (
  .O(mux_o_170),
  .I0(dpx9b_inst_20_douta[24]),
  .I1(dpx9b_inst_21_douta[24]),
  .S0(dff_q_2)
);
MUX2 mux_inst_171 (
  .O(mux_o_171),
  .I0(dpx9b_inst_22_douta[24]),
  .I1(dpx9b_inst_23_douta[24]),
  .S0(dff_q_2)
);
MUX2 mux_inst_172 (
  .O(mux_o_172),
  .I0(mux_o_168),
  .I1(mux_o_169),
  .S0(dff_q_1)
);
MUX2 mux_inst_173 (
  .O(mux_o_173),
  .I0(mux_o_170),
  .I1(mux_o_171),
  .S0(dff_q_1)
);
MUX2 mux_inst_174 (
  .O(douta[24]),
  .I0(mux_o_172),
  .I1(mux_o_173),
  .S0(dff_q_0)
);
MUX2 mux_inst_175 (
  .O(mux_o_175),
  .I0(dpx9b_inst_16_douta[25]),
  .I1(dpx9b_inst_17_douta[25]),
  .S0(dff_q_2)
);
MUX2 mux_inst_176 (
  .O(mux_o_176),
  .I0(dpx9b_inst_18_douta[25]),
  .I1(dpx9b_inst_19_douta[25]),
  .S0(dff_q_2)
);
MUX2 mux_inst_177 (
  .O(mux_o_177),
  .I0(dpx9b_inst_20_douta[25]),
  .I1(dpx9b_inst_21_douta[25]),
  .S0(dff_q_2)
);
MUX2 mux_inst_178 (
  .O(mux_o_178),
  .I0(dpx9b_inst_22_douta[25]),
  .I1(dpx9b_inst_23_douta[25]),
  .S0(dff_q_2)
);
MUX2 mux_inst_179 (
  .O(mux_o_179),
  .I0(mux_o_175),
  .I1(mux_o_176),
  .S0(dff_q_1)
);
MUX2 mux_inst_180 (
  .O(mux_o_180),
  .I0(mux_o_177),
  .I1(mux_o_178),
  .S0(dff_q_1)
);
MUX2 mux_inst_181 (
  .O(douta[25]),
  .I0(mux_o_179),
  .I1(mux_o_180),
  .S0(dff_q_0)
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(dpx9b_inst_16_douta[26]),
  .I1(dpx9b_inst_17_douta[26]),
  .S0(dff_q_2)
);
MUX2 mux_inst_183 (
  .O(mux_o_183),
  .I0(dpx9b_inst_18_douta[26]),
  .I1(dpx9b_inst_19_douta[26]),
  .S0(dff_q_2)
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(dpx9b_inst_20_douta[26]),
  .I1(dpx9b_inst_21_douta[26]),
  .S0(dff_q_2)
);
MUX2 mux_inst_185 (
  .O(mux_o_185),
  .I0(dpx9b_inst_22_douta[26]),
  .I1(dpx9b_inst_23_douta[26]),
  .S0(dff_q_2)
);
MUX2 mux_inst_186 (
  .O(mux_o_186),
  .I0(mux_o_182),
  .I1(mux_o_183),
  .S0(dff_q_1)
);
MUX2 mux_inst_187 (
  .O(mux_o_187),
  .I0(mux_o_184),
  .I1(mux_o_185),
  .S0(dff_q_1)
);
MUX2 mux_inst_188 (
  .O(douta[26]),
  .I0(mux_o_186),
  .I1(mux_o_187),
  .S0(dff_q_0)
);
MUX2 mux_inst_189 (
  .O(mux_o_189),
  .I0(dpx9b_inst_0_doutb[0]),
  .I1(dpx9b_inst_1_doutb[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_190 (
  .O(mux_o_190),
  .I0(dpx9b_inst_2_doutb[0]),
  .I1(dpx9b_inst_3_doutb[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_191 (
  .O(mux_o_191),
  .I0(dpx9b_inst_4_doutb[0]),
  .I1(dpx9b_inst_5_doutb[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_192 (
  .O(mux_o_192),
  .I0(dpx9b_inst_6_doutb[0]),
  .I1(dpx9b_inst_7_doutb[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_193 (
  .O(mux_o_193),
  .I0(mux_o_189),
  .I1(mux_o_190),
  .S0(dff_q_4)
);
MUX2 mux_inst_194 (
  .O(mux_o_194),
  .I0(mux_o_191),
  .I1(mux_o_192),
  .S0(dff_q_4)
);
MUX2 mux_inst_195 (
  .O(doutb[0]),
  .I0(mux_o_193),
  .I1(mux_o_194),
  .S0(dff_q_3)
);
MUX2 mux_inst_196 (
  .O(mux_o_196),
  .I0(dpx9b_inst_0_doutb[1]),
  .I1(dpx9b_inst_1_doutb[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_197 (
  .O(mux_o_197),
  .I0(dpx9b_inst_2_doutb[1]),
  .I1(dpx9b_inst_3_doutb[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_198 (
  .O(mux_o_198),
  .I0(dpx9b_inst_4_doutb[1]),
  .I1(dpx9b_inst_5_doutb[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_199 (
  .O(mux_o_199),
  .I0(dpx9b_inst_6_doutb[1]),
  .I1(dpx9b_inst_7_doutb[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_200 (
  .O(mux_o_200),
  .I0(mux_o_196),
  .I1(mux_o_197),
  .S0(dff_q_4)
);
MUX2 mux_inst_201 (
  .O(mux_o_201),
  .I0(mux_o_198),
  .I1(mux_o_199),
  .S0(dff_q_4)
);
MUX2 mux_inst_202 (
  .O(doutb[1]),
  .I0(mux_o_200),
  .I1(mux_o_201),
  .S0(dff_q_3)
);
MUX2 mux_inst_203 (
  .O(mux_o_203),
  .I0(dpx9b_inst_0_doutb[2]),
  .I1(dpx9b_inst_1_doutb[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_204 (
  .O(mux_o_204),
  .I0(dpx9b_inst_2_doutb[2]),
  .I1(dpx9b_inst_3_doutb[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_205 (
  .O(mux_o_205),
  .I0(dpx9b_inst_4_doutb[2]),
  .I1(dpx9b_inst_5_doutb[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_206 (
  .O(mux_o_206),
  .I0(dpx9b_inst_6_doutb[2]),
  .I1(dpx9b_inst_7_doutb[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_207 (
  .O(mux_o_207),
  .I0(mux_o_203),
  .I1(mux_o_204),
  .S0(dff_q_4)
);
MUX2 mux_inst_208 (
  .O(mux_o_208),
  .I0(mux_o_205),
  .I1(mux_o_206),
  .S0(dff_q_4)
);
MUX2 mux_inst_209 (
  .O(doutb[2]),
  .I0(mux_o_207),
  .I1(mux_o_208),
  .S0(dff_q_3)
);
MUX2 mux_inst_210 (
  .O(mux_o_210),
  .I0(dpx9b_inst_0_doutb[3]),
  .I1(dpx9b_inst_1_doutb[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_211 (
  .O(mux_o_211),
  .I0(dpx9b_inst_2_doutb[3]),
  .I1(dpx9b_inst_3_doutb[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_212 (
  .O(mux_o_212),
  .I0(dpx9b_inst_4_doutb[3]),
  .I1(dpx9b_inst_5_doutb[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_213 (
  .O(mux_o_213),
  .I0(dpx9b_inst_6_doutb[3]),
  .I1(dpx9b_inst_7_doutb[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_214 (
  .O(mux_o_214),
  .I0(mux_o_210),
  .I1(mux_o_211),
  .S0(dff_q_4)
);
MUX2 mux_inst_215 (
  .O(mux_o_215),
  .I0(mux_o_212),
  .I1(mux_o_213),
  .S0(dff_q_4)
);
MUX2 mux_inst_216 (
  .O(doutb[3]),
  .I0(mux_o_214),
  .I1(mux_o_215),
  .S0(dff_q_3)
);
MUX2 mux_inst_217 (
  .O(mux_o_217),
  .I0(dpx9b_inst_0_doutb[4]),
  .I1(dpx9b_inst_1_doutb[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_218 (
  .O(mux_o_218),
  .I0(dpx9b_inst_2_doutb[4]),
  .I1(dpx9b_inst_3_doutb[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_219 (
  .O(mux_o_219),
  .I0(dpx9b_inst_4_doutb[4]),
  .I1(dpx9b_inst_5_doutb[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_220 (
  .O(mux_o_220),
  .I0(dpx9b_inst_6_doutb[4]),
  .I1(dpx9b_inst_7_doutb[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_221 (
  .O(mux_o_221),
  .I0(mux_o_217),
  .I1(mux_o_218),
  .S0(dff_q_4)
);
MUX2 mux_inst_222 (
  .O(mux_o_222),
  .I0(mux_o_219),
  .I1(mux_o_220),
  .S0(dff_q_4)
);
MUX2 mux_inst_223 (
  .O(doutb[4]),
  .I0(mux_o_221),
  .I1(mux_o_222),
  .S0(dff_q_3)
);
MUX2 mux_inst_224 (
  .O(mux_o_224),
  .I0(dpx9b_inst_0_doutb[5]),
  .I1(dpx9b_inst_1_doutb[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_225 (
  .O(mux_o_225),
  .I0(dpx9b_inst_2_doutb[5]),
  .I1(dpx9b_inst_3_doutb[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_226 (
  .O(mux_o_226),
  .I0(dpx9b_inst_4_doutb[5]),
  .I1(dpx9b_inst_5_doutb[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_227 (
  .O(mux_o_227),
  .I0(dpx9b_inst_6_doutb[5]),
  .I1(dpx9b_inst_7_doutb[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_228 (
  .O(mux_o_228),
  .I0(mux_o_224),
  .I1(mux_o_225),
  .S0(dff_q_4)
);
MUX2 mux_inst_229 (
  .O(mux_o_229),
  .I0(mux_o_226),
  .I1(mux_o_227),
  .S0(dff_q_4)
);
MUX2 mux_inst_230 (
  .O(doutb[5]),
  .I0(mux_o_228),
  .I1(mux_o_229),
  .S0(dff_q_3)
);
MUX2 mux_inst_231 (
  .O(mux_o_231),
  .I0(dpx9b_inst_0_doutb[6]),
  .I1(dpx9b_inst_1_doutb[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_232 (
  .O(mux_o_232),
  .I0(dpx9b_inst_2_doutb[6]),
  .I1(dpx9b_inst_3_doutb[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_233 (
  .O(mux_o_233),
  .I0(dpx9b_inst_4_doutb[6]),
  .I1(dpx9b_inst_5_doutb[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_234 (
  .O(mux_o_234),
  .I0(dpx9b_inst_6_doutb[6]),
  .I1(dpx9b_inst_7_doutb[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_235 (
  .O(mux_o_235),
  .I0(mux_o_231),
  .I1(mux_o_232),
  .S0(dff_q_4)
);
MUX2 mux_inst_236 (
  .O(mux_o_236),
  .I0(mux_o_233),
  .I1(mux_o_234),
  .S0(dff_q_4)
);
MUX2 mux_inst_237 (
  .O(doutb[6]),
  .I0(mux_o_235),
  .I1(mux_o_236),
  .S0(dff_q_3)
);
MUX2 mux_inst_238 (
  .O(mux_o_238),
  .I0(dpx9b_inst_0_doutb[7]),
  .I1(dpx9b_inst_1_doutb[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_239 (
  .O(mux_o_239),
  .I0(dpx9b_inst_2_doutb[7]),
  .I1(dpx9b_inst_3_doutb[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_240 (
  .O(mux_o_240),
  .I0(dpx9b_inst_4_doutb[7]),
  .I1(dpx9b_inst_5_doutb[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_241 (
  .O(mux_o_241),
  .I0(dpx9b_inst_6_doutb[7]),
  .I1(dpx9b_inst_7_doutb[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_242 (
  .O(mux_o_242),
  .I0(mux_o_238),
  .I1(mux_o_239),
  .S0(dff_q_4)
);
MUX2 mux_inst_243 (
  .O(mux_o_243),
  .I0(mux_o_240),
  .I1(mux_o_241),
  .S0(dff_q_4)
);
MUX2 mux_inst_244 (
  .O(doutb[7]),
  .I0(mux_o_242),
  .I1(mux_o_243),
  .S0(dff_q_3)
);
MUX2 mux_inst_245 (
  .O(mux_o_245),
  .I0(dpx9b_inst_0_doutb[8]),
  .I1(dpx9b_inst_1_doutb[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_246 (
  .O(mux_o_246),
  .I0(dpx9b_inst_2_doutb[8]),
  .I1(dpx9b_inst_3_doutb[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_247 (
  .O(mux_o_247),
  .I0(dpx9b_inst_4_doutb[8]),
  .I1(dpx9b_inst_5_doutb[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_248 (
  .O(mux_o_248),
  .I0(dpx9b_inst_6_doutb[8]),
  .I1(dpx9b_inst_7_doutb[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_249 (
  .O(mux_o_249),
  .I0(mux_o_245),
  .I1(mux_o_246),
  .S0(dff_q_4)
);
MUX2 mux_inst_250 (
  .O(mux_o_250),
  .I0(mux_o_247),
  .I1(mux_o_248),
  .S0(dff_q_4)
);
MUX2 mux_inst_251 (
  .O(doutb[8]),
  .I0(mux_o_249),
  .I1(mux_o_250),
  .S0(dff_q_3)
);
MUX2 mux_inst_252 (
  .O(mux_o_252),
  .I0(dpx9b_inst_8_doutb[9]),
  .I1(dpx9b_inst_9_doutb[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_253 (
  .O(mux_o_253),
  .I0(dpx9b_inst_10_doutb[9]),
  .I1(dpx9b_inst_11_doutb[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_254 (
  .O(mux_o_254),
  .I0(dpx9b_inst_12_doutb[9]),
  .I1(dpx9b_inst_13_doutb[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_255 (
  .O(mux_o_255),
  .I0(dpx9b_inst_14_doutb[9]),
  .I1(dpx9b_inst_15_doutb[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_256 (
  .O(mux_o_256),
  .I0(mux_o_252),
  .I1(mux_o_253),
  .S0(dff_q_4)
);
MUX2 mux_inst_257 (
  .O(mux_o_257),
  .I0(mux_o_254),
  .I1(mux_o_255),
  .S0(dff_q_4)
);
MUX2 mux_inst_258 (
  .O(doutb[9]),
  .I0(mux_o_256),
  .I1(mux_o_257),
  .S0(dff_q_3)
);
MUX2 mux_inst_259 (
  .O(mux_o_259),
  .I0(dpx9b_inst_8_doutb[10]),
  .I1(dpx9b_inst_9_doutb[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_260 (
  .O(mux_o_260),
  .I0(dpx9b_inst_10_doutb[10]),
  .I1(dpx9b_inst_11_doutb[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_261 (
  .O(mux_o_261),
  .I0(dpx9b_inst_12_doutb[10]),
  .I1(dpx9b_inst_13_doutb[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_262 (
  .O(mux_o_262),
  .I0(dpx9b_inst_14_doutb[10]),
  .I1(dpx9b_inst_15_doutb[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_263 (
  .O(mux_o_263),
  .I0(mux_o_259),
  .I1(mux_o_260),
  .S0(dff_q_4)
);
MUX2 mux_inst_264 (
  .O(mux_o_264),
  .I0(mux_o_261),
  .I1(mux_o_262),
  .S0(dff_q_4)
);
MUX2 mux_inst_265 (
  .O(doutb[10]),
  .I0(mux_o_263),
  .I1(mux_o_264),
  .S0(dff_q_3)
);
MUX2 mux_inst_266 (
  .O(mux_o_266),
  .I0(dpx9b_inst_8_doutb[11]),
  .I1(dpx9b_inst_9_doutb[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_267 (
  .O(mux_o_267),
  .I0(dpx9b_inst_10_doutb[11]),
  .I1(dpx9b_inst_11_doutb[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_268 (
  .O(mux_o_268),
  .I0(dpx9b_inst_12_doutb[11]),
  .I1(dpx9b_inst_13_doutb[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_269 (
  .O(mux_o_269),
  .I0(dpx9b_inst_14_doutb[11]),
  .I1(dpx9b_inst_15_doutb[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_270 (
  .O(mux_o_270),
  .I0(mux_o_266),
  .I1(mux_o_267),
  .S0(dff_q_4)
);
MUX2 mux_inst_271 (
  .O(mux_o_271),
  .I0(mux_o_268),
  .I1(mux_o_269),
  .S0(dff_q_4)
);
MUX2 mux_inst_272 (
  .O(doutb[11]),
  .I0(mux_o_270),
  .I1(mux_o_271),
  .S0(dff_q_3)
);
MUX2 mux_inst_273 (
  .O(mux_o_273),
  .I0(dpx9b_inst_8_doutb[12]),
  .I1(dpx9b_inst_9_doutb[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_274 (
  .O(mux_o_274),
  .I0(dpx9b_inst_10_doutb[12]),
  .I1(dpx9b_inst_11_doutb[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_275 (
  .O(mux_o_275),
  .I0(dpx9b_inst_12_doutb[12]),
  .I1(dpx9b_inst_13_doutb[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_276 (
  .O(mux_o_276),
  .I0(dpx9b_inst_14_doutb[12]),
  .I1(dpx9b_inst_15_doutb[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_277 (
  .O(mux_o_277),
  .I0(mux_o_273),
  .I1(mux_o_274),
  .S0(dff_q_4)
);
MUX2 mux_inst_278 (
  .O(mux_o_278),
  .I0(mux_o_275),
  .I1(mux_o_276),
  .S0(dff_q_4)
);
MUX2 mux_inst_279 (
  .O(doutb[12]),
  .I0(mux_o_277),
  .I1(mux_o_278),
  .S0(dff_q_3)
);
MUX2 mux_inst_280 (
  .O(mux_o_280),
  .I0(dpx9b_inst_8_doutb[13]),
  .I1(dpx9b_inst_9_doutb[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_281 (
  .O(mux_o_281),
  .I0(dpx9b_inst_10_doutb[13]),
  .I1(dpx9b_inst_11_doutb[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_282 (
  .O(mux_o_282),
  .I0(dpx9b_inst_12_doutb[13]),
  .I1(dpx9b_inst_13_doutb[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_283 (
  .O(mux_o_283),
  .I0(dpx9b_inst_14_doutb[13]),
  .I1(dpx9b_inst_15_doutb[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_284 (
  .O(mux_o_284),
  .I0(mux_o_280),
  .I1(mux_o_281),
  .S0(dff_q_4)
);
MUX2 mux_inst_285 (
  .O(mux_o_285),
  .I0(mux_o_282),
  .I1(mux_o_283),
  .S0(dff_q_4)
);
MUX2 mux_inst_286 (
  .O(doutb[13]),
  .I0(mux_o_284),
  .I1(mux_o_285),
  .S0(dff_q_3)
);
MUX2 mux_inst_287 (
  .O(mux_o_287),
  .I0(dpx9b_inst_8_doutb[14]),
  .I1(dpx9b_inst_9_doutb[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_288 (
  .O(mux_o_288),
  .I0(dpx9b_inst_10_doutb[14]),
  .I1(dpx9b_inst_11_doutb[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_289 (
  .O(mux_o_289),
  .I0(dpx9b_inst_12_doutb[14]),
  .I1(dpx9b_inst_13_doutb[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_290 (
  .O(mux_o_290),
  .I0(dpx9b_inst_14_doutb[14]),
  .I1(dpx9b_inst_15_doutb[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_291 (
  .O(mux_o_291),
  .I0(mux_o_287),
  .I1(mux_o_288),
  .S0(dff_q_4)
);
MUX2 mux_inst_292 (
  .O(mux_o_292),
  .I0(mux_o_289),
  .I1(mux_o_290),
  .S0(dff_q_4)
);
MUX2 mux_inst_293 (
  .O(doutb[14]),
  .I0(mux_o_291),
  .I1(mux_o_292),
  .S0(dff_q_3)
);
MUX2 mux_inst_294 (
  .O(mux_o_294),
  .I0(dpx9b_inst_8_doutb[15]),
  .I1(dpx9b_inst_9_doutb[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_295 (
  .O(mux_o_295),
  .I0(dpx9b_inst_10_doutb[15]),
  .I1(dpx9b_inst_11_doutb[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_296 (
  .O(mux_o_296),
  .I0(dpx9b_inst_12_doutb[15]),
  .I1(dpx9b_inst_13_doutb[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_297 (
  .O(mux_o_297),
  .I0(dpx9b_inst_14_doutb[15]),
  .I1(dpx9b_inst_15_doutb[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_298 (
  .O(mux_o_298),
  .I0(mux_o_294),
  .I1(mux_o_295),
  .S0(dff_q_4)
);
MUX2 mux_inst_299 (
  .O(mux_o_299),
  .I0(mux_o_296),
  .I1(mux_o_297),
  .S0(dff_q_4)
);
MUX2 mux_inst_300 (
  .O(doutb[15]),
  .I0(mux_o_298),
  .I1(mux_o_299),
  .S0(dff_q_3)
);
MUX2 mux_inst_301 (
  .O(mux_o_301),
  .I0(dpx9b_inst_8_doutb[16]),
  .I1(dpx9b_inst_9_doutb[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_302 (
  .O(mux_o_302),
  .I0(dpx9b_inst_10_doutb[16]),
  .I1(dpx9b_inst_11_doutb[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_303 (
  .O(mux_o_303),
  .I0(dpx9b_inst_12_doutb[16]),
  .I1(dpx9b_inst_13_doutb[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_304 (
  .O(mux_o_304),
  .I0(dpx9b_inst_14_doutb[16]),
  .I1(dpx9b_inst_15_doutb[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_305 (
  .O(mux_o_305),
  .I0(mux_o_301),
  .I1(mux_o_302),
  .S0(dff_q_4)
);
MUX2 mux_inst_306 (
  .O(mux_o_306),
  .I0(mux_o_303),
  .I1(mux_o_304),
  .S0(dff_q_4)
);
MUX2 mux_inst_307 (
  .O(doutb[16]),
  .I0(mux_o_305),
  .I1(mux_o_306),
  .S0(dff_q_3)
);
MUX2 mux_inst_308 (
  .O(mux_o_308),
  .I0(dpx9b_inst_8_doutb[17]),
  .I1(dpx9b_inst_9_doutb[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_309 (
  .O(mux_o_309),
  .I0(dpx9b_inst_10_doutb[17]),
  .I1(dpx9b_inst_11_doutb[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_310 (
  .O(mux_o_310),
  .I0(dpx9b_inst_12_doutb[17]),
  .I1(dpx9b_inst_13_doutb[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_311 (
  .O(mux_o_311),
  .I0(dpx9b_inst_14_doutb[17]),
  .I1(dpx9b_inst_15_doutb[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_312 (
  .O(mux_o_312),
  .I0(mux_o_308),
  .I1(mux_o_309),
  .S0(dff_q_4)
);
MUX2 mux_inst_313 (
  .O(mux_o_313),
  .I0(mux_o_310),
  .I1(mux_o_311),
  .S0(dff_q_4)
);
MUX2 mux_inst_314 (
  .O(doutb[17]),
  .I0(mux_o_312),
  .I1(mux_o_313),
  .S0(dff_q_3)
);
MUX2 mux_inst_315 (
  .O(mux_o_315),
  .I0(dpx9b_inst_16_doutb[18]),
  .I1(dpx9b_inst_17_doutb[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_316 (
  .O(mux_o_316),
  .I0(dpx9b_inst_18_doutb[18]),
  .I1(dpx9b_inst_19_doutb[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_317 (
  .O(mux_o_317),
  .I0(dpx9b_inst_20_doutb[18]),
  .I1(dpx9b_inst_21_doutb[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_318 (
  .O(mux_o_318),
  .I0(dpx9b_inst_22_doutb[18]),
  .I1(dpx9b_inst_23_doutb[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_319 (
  .O(mux_o_319),
  .I0(mux_o_315),
  .I1(mux_o_316),
  .S0(dff_q_4)
);
MUX2 mux_inst_320 (
  .O(mux_o_320),
  .I0(mux_o_317),
  .I1(mux_o_318),
  .S0(dff_q_4)
);
MUX2 mux_inst_321 (
  .O(doutb[18]),
  .I0(mux_o_319),
  .I1(mux_o_320),
  .S0(dff_q_3)
);
MUX2 mux_inst_322 (
  .O(mux_o_322),
  .I0(dpx9b_inst_16_doutb[19]),
  .I1(dpx9b_inst_17_doutb[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_323 (
  .O(mux_o_323),
  .I0(dpx9b_inst_18_doutb[19]),
  .I1(dpx9b_inst_19_doutb[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_324 (
  .O(mux_o_324),
  .I0(dpx9b_inst_20_doutb[19]),
  .I1(dpx9b_inst_21_doutb[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_325 (
  .O(mux_o_325),
  .I0(dpx9b_inst_22_doutb[19]),
  .I1(dpx9b_inst_23_doutb[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_326 (
  .O(mux_o_326),
  .I0(mux_o_322),
  .I1(mux_o_323),
  .S0(dff_q_4)
);
MUX2 mux_inst_327 (
  .O(mux_o_327),
  .I0(mux_o_324),
  .I1(mux_o_325),
  .S0(dff_q_4)
);
MUX2 mux_inst_328 (
  .O(doutb[19]),
  .I0(mux_o_326),
  .I1(mux_o_327),
  .S0(dff_q_3)
);
MUX2 mux_inst_329 (
  .O(mux_o_329),
  .I0(dpx9b_inst_16_doutb[20]),
  .I1(dpx9b_inst_17_doutb[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_330 (
  .O(mux_o_330),
  .I0(dpx9b_inst_18_doutb[20]),
  .I1(dpx9b_inst_19_doutb[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_331 (
  .O(mux_o_331),
  .I0(dpx9b_inst_20_doutb[20]),
  .I1(dpx9b_inst_21_doutb[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_332 (
  .O(mux_o_332),
  .I0(dpx9b_inst_22_doutb[20]),
  .I1(dpx9b_inst_23_doutb[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_333 (
  .O(mux_o_333),
  .I0(mux_o_329),
  .I1(mux_o_330),
  .S0(dff_q_4)
);
MUX2 mux_inst_334 (
  .O(mux_o_334),
  .I0(mux_o_331),
  .I1(mux_o_332),
  .S0(dff_q_4)
);
MUX2 mux_inst_335 (
  .O(doutb[20]),
  .I0(mux_o_333),
  .I1(mux_o_334),
  .S0(dff_q_3)
);
MUX2 mux_inst_336 (
  .O(mux_o_336),
  .I0(dpx9b_inst_16_doutb[21]),
  .I1(dpx9b_inst_17_doutb[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_337 (
  .O(mux_o_337),
  .I0(dpx9b_inst_18_doutb[21]),
  .I1(dpx9b_inst_19_doutb[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_338 (
  .O(mux_o_338),
  .I0(dpx9b_inst_20_doutb[21]),
  .I1(dpx9b_inst_21_doutb[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_339 (
  .O(mux_o_339),
  .I0(dpx9b_inst_22_doutb[21]),
  .I1(dpx9b_inst_23_doutb[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_340 (
  .O(mux_o_340),
  .I0(mux_o_336),
  .I1(mux_o_337),
  .S0(dff_q_4)
);
MUX2 mux_inst_341 (
  .O(mux_o_341),
  .I0(mux_o_338),
  .I1(mux_o_339),
  .S0(dff_q_4)
);
MUX2 mux_inst_342 (
  .O(doutb[21]),
  .I0(mux_o_340),
  .I1(mux_o_341),
  .S0(dff_q_3)
);
MUX2 mux_inst_343 (
  .O(mux_o_343),
  .I0(dpx9b_inst_16_doutb[22]),
  .I1(dpx9b_inst_17_doutb[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_344 (
  .O(mux_o_344),
  .I0(dpx9b_inst_18_doutb[22]),
  .I1(dpx9b_inst_19_doutb[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_345 (
  .O(mux_o_345),
  .I0(dpx9b_inst_20_doutb[22]),
  .I1(dpx9b_inst_21_doutb[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_346 (
  .O(mux_o_346),
  .I0(dpx9b_inst_22_doutb[22]),
  .I1(dpx9b_inst_23_doutb[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_347 (
  .O(mux_o_347),
  .I0(mux_o_343),
  .I1(mux_o_344),
  .S0(dff_q_4)
);
MUX2 mux_inst_348 (
  .O(mux_o_348),
  .I0(mux_o_345),
  .I1(mux_o_346),
  .S0(dff_q_4)
);
MUX2 mux_inst_349 (
  .O(doutb[22]),
  .I0(mux_o_347),
  .I1(mux_o_348),
  .S0(dff_q_3)
);
MUX2 mux_inst_350 (
  .O(mux_o_350),
  .I0(dpx9b_inst_16_doutb[23]),
  .I1(dpx9b_inst_17_doutb[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_351 (
  .O(mux_o_351),
  .I0(dpx9b_inst_18_doutb[23]),
  .I1(dpx9b_inst_19_doutb[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_352 (
  .O(mux_o_352),
  .I0(dpx9b_inst_20_doutb[23]),
  .I1(dpx9b_inst_21_doutb[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_353 (
  .O(mux_o_353),
  .I0(dpx9b_inst_22_doutb[23]),
  .I1(dpx9b_inst_23_doutb[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_354 (
  .O(mux_o_354),
  .I0(mux_o_350),
  .I1(mux_o_351),
  .S0(dff_q_4)
);
MUX2 mux_inst_355 (
  .O(mux_o_355),
  .I0(mux_o_352),
  .I1(mux_o_353),
  .S0(dff_q_4)
);
MUX2 mux_inst_356 (
  .O(doutb[23]),
  .I0(mux_o_354),
  .I1(mux_o_355),
  .S0(dff_q_3)
);
MUX2 mux_inst_357 (
  .O(mux_o_357),
  .I0(dpx9b_inst_16_doutb[24]),
  .I1(dpx9b_inst_17_doutb[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_358 (
  .O(mux_o_358),
  .I0(dpx9b_inst_18_doutb[24]),
  .I1(dpx9b_inst_19_doutb[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_359 (
  .O(mux_o_359),
  .I0(dpx9b_inst_20_doutb[24]),
  .I1(dpx9b_inst_21_doutb[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_360 (
  .O(mux_o_360),
  .I0(dpx9b_inst_22_doutb[24]),
  .I1(dpx9b_inst_23_doutb[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_361 (
  .O(mux_o_361),
  .I0(mux_o_357),
  .I1(mux_o_358),
  .S0(dff_q_4)
);
MUX2 mux_inst_362 (
  .O(mux_o_362),
  .I0(mux_o_359),
  .I1(mux_o_360),
  .S0(dff_q_4)
);
MUX2 mux_inst_363 (
  .O(doutb[24]),
  .I0(mux_o_361),
  .I1(mux_o_362),
  .S0(dff_q_3)
);
MUX2 mux_inst_364 (
  .O(mux_o_364),
  .I0(dpx9b_inst_16_doutb[25]),
  .I1(dpx9b_inst_17_doutb[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_365 (
  .O(mux_o_365),
  .I0(dpx9b_inst_18_doutb[25]),
  .I1(dpx9b_inst_19_doutb[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_366 (
  .O(mux_o_366),
  .I0(dpx9b_inst_20_doutb[25]),
  .I1(dpx9b_inst_21_doutb[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_367 (
  .O(mux_o_367),
  .I0(dpx9b_inst_22_doutb[25]),
  .I1(dpx9b_inst_23_doutb[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_368 (
  .O(mux_o_368),
  .I0(mux_o_364),
  .I1(mux_o_365),
  .S0(dff_q_4)
);
MUX2 mux_inst_369 (
  .O(mux_o_369),
  .I0(mux_o_366),
  .I1(mux_o_367),
  .S0(dff_q_4)
);
MUX2 mux_inst_370 (
  .O(doutb[25]),
  .I0(mux_o_368),
  .I1(mux_o_369),
  .S0(dff_q_3)
);
MUX2 mux_inst_371 (
  .O(mux_o_371),
  .I0(dpx9b_inst_16_doutb[26]),
  .I1(dpx9b_inst_17_doutb[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_372 (
  .O(mux_o_372),
  .I0(dpx9b_inst_18_doutb[26]),
  .I1(dpx9b_inst_19_doutb[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_373 (
  .O(mux_o_373),
  .I0(dpx9b_inst_20_doutb[26]),
  .I1(dpx9b_inst_21_doutb[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_374 (
  .O(mux_o_374),
  .I0(dpx9b_inst_22_doutb[26]),
  .I1(dpx9b_inst_23_doutb[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_375 (
  .O(mux_o_375),
  .I0(mux_o_371),
  .I1(mux_o_372),
  .S0(dff_q_4)
);
MUX2 mux_inst_376 (
  .O(mux_o_376),
  .I0(mux_o_373),
  .I1(mux_o_374),
  .S0(dff_q_4)
);
MUX2 mux_inst_377 (
  .O(doutb[26]),
  .I0(mux_o_375),
  .I1(mux_o_376),
  .S0(dff_q_3)
);
endmodule //Gowin_DPB
