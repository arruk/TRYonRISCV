TORVS/torvs1.sv