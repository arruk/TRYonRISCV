module adder8b(
	input[7:0] a,
	input[7:0] b,
	output [7:0] s,
	output cout
);



endmodule
