TORVS/core.sv